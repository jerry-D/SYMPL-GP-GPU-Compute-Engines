-- Copyright 2003-2006 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package pkg_fp_exp_exp_y2 is

  component fp_exp_exp_y2_6 is
    port ( nY2    : in  std_logic_vector(2 downto 0);
           nExpY2 : out std_logic_vector(2 downto 0) );
  end component;

  component fp_exp_exp_y2_7 is
    port ( nY2    : in  std_logic_vector(3 downto 0);
           nExpY2 : out std_logic_vector(3 downto 0) );
  end component;

  component fp_exp_exp_y2_8 is
    port ( nY2    : in  std_logic_vector(4 downto 0);
           nExpY2 : out std_logic_vector(4 downto 0) );
  end component;

  component fp_exp_exp_y2_9 is
    port ( nY2    : in  std_logic_vector(3 downto 0);
           nExpY2 : out std_logic_vector(3 downto 0) );
  end component;

  component fp_exp_exp_y2_10 is
    port ( nY2    : in  std_logic_vector(4 downto 0);
           nExpY2 : out std_logic_vector(4 downto 0) );
  end component;

  component fp_exp_exp_y2_11 is
    port ( nY2    : in  std_logic_vector(5 downto 0);
           nExpY2 : out std_logic_vector(5 downto 0) );
  end component;

  component fp_exp_exp_y2_12 is
    port ( nY2    : in  std_logic_vector(4 downto 0);
           nExpY2 : out std_logic_vector(4 downto 0) );
  end component;

  component fp_exp_exp_y2_13 is
    port ( nY2    : in  std_logic_vector(5 downto 0);
           nExpY2 : out std_logic_vector(5 downto 0) );
  end component;

  component fp_exp_exp_y2_14 is
    port ( nY2    : in  std_logic_vector(6 downto 0);
           nExpY2 : out std_logic_vector(6 downto 0) );
  end component;

  component fp_exp_exp_y2_15 is
    port ( nY2    : in  std_logic_vector(5 downto 0);
           nExpY2 : out std_logic_vector(5 downto 0) );
  end component;

  component fp_exp_exp_y2_16 is
    port ( nY2    : in  std_logic_vector(6 downto 0);
           nExpY2 : out std_logic_vector(6 downto 0) );
  end component;

  component fp_exp_exp_y2_17 is
    port ( nY2    : in  std_logic_vector(7 downto 0);
           nExpY2 : out std_logic_vector(7 downto 0) );
  end component;

  component fp_exp_exp_y2_18 is
    port ( nY2    : in  std_logic_vector(6 downto 0);
           nExpY2 : out std_logic_vector(6 downto 0) );
  end component;

  component fp_exp_exp_y2_19 is
    port ( nY2    : in  std_logic_vector(7 downto 0);
           nExpY2 : out std_logic_vector(7 downto 0) );
  end component;

  component fp_exp_exp_y2_20 is
    port ( x : in  std_logic_vector(8 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component fp_exp_exp_y2_20_clk is
    port ( x   : in  std_logic_vector(8 downto 0);
           r   : out std_logic_vector(9 downto 0);
           clk : in  std_logic );
  end component;

  component fp_exp_exp_y2_21 is
    port ( x : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component fp_exp_exp_y2_21_clk is
    port ( x   : in  std_logic_vector(9 downto 0);
           r   : out std_logic_vector(10 downto 0);
           clk : in  std_logic );
  end component;

  component fp_exp_exp_y2_22 is
    port ( x : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component fp_exp_exp_y2_22_clk is
    port ( x   : in  std_logic_vector(10 downto 0);
           r   : out std_logic_vector(11 downto 0);
           clk : in  std_logic );
  end component;

  component fp_exp_exp_y2_23 is
    port ( x : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  component fp_exp_exp_y2_23_clk is
    port ( x   : in  std_logic_vector(11 downto 0);
           r   : out std_logic_vector(12 downto 0);
           clk : in  std_logic );
  end component;

end package;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_6 is
  port ( nY2    : in  std_logic_vector(2 downto 0);
         nExpY2 : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_6 is
begin

  with nY2 select
    nExpY2 <= "000" when "000", -- t[0] = 0
              "000" when "001", -- t[1] = 0
              "000" when "010", -- t[2] = 0
              "001" when "011", -- t[3] = 1
              "001" when "100", -- t[4] = 1
              "010" when "101", -- t[5] = 2
              "010" when "110", -- t[6] = 2
              "011" when "111", -- t[7] = 3
              "---" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_7 is
  port ( nY2    : in  std_logic_vector(3 downto 0);
         nExpY2 : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_7 is
begin

  with nY2 select
    nExpY2 <= "0000" when "0000", -- t[0] = 0
              "0000" when "0001", -- t[1] = 0
              "0000" when "0010", -- t[2] = 0
              "0000" when "0011", -- t[3] = 0
              "0001" when "0100", -- t[4] = 1
              "0001" when "0101", -- t[5] = 1
              "0001" when "0110", -- t[6] = 1
              "0010" when "0111", -- t[7] = 2
              "0010" when "1000", -- t[8] = 2
              "0011" when "1001", -- t[9] = 3
              "0011" when "1010", -- t[10] = 3
              "0100" when "1011", -- t[11] = 4
              "0101" when "1100", -- t[12] = 5
              "0101" when "1101", -- t[13] = 5
              "0110" when "1110", -- t[14] = 6
              "0111" when "1111", -- t[15] = 7
              "----" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_8 is
  port ( nY2    : in  std_logic_vector(4 downto 0);
         nExpY2 : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_8 is
begin

  with nY2 select
    nExpY2 <= "00000" when "00000", -- t[0] = 0
              "00000" when "00001", -- t[1] = 0
              "00000" when "00010", -- t[2] = 0
              "00000" when "00011", -- t[3] = 0
              "00000" when "00100", -- t[4] = 0
              "00000" when "00101", -- t[5] = 0
              "00001" when "00110", -- t[6] = 1
              "00001" when "00111", -- t[7] = 1
              "00001" when "01000", -- t[8] = 1
              "00001" when "01001", -- t[9] = 1
              "00010" when "01010", -- t[10] = 2
              "00010" when "01011", -- t[11] = 2
              "00010" when "01100", -- t[12] = 2
              "00011" when "01101", -- t[13] = 3
              "00011" when "01110", -- t[14] = 3
              "00100" when "01111", -- t[15] = 4
              "00100" when "10000", -- t[16] = 4
              "00101" when "10001", -- t[17] = 5
              "00101" when "10010", -- t[18] = 5
              "00110" when "10011", -- t[19] = 6
              "00110" when "10100", -- t[20] = 6
              "00111" when "10101", -- t[21] = 7
              "01000" when "10110", -- t[22] = 8
              "01000" when "10111", -- t[23] = 8
              "01001" when "11000", -- t[24] = 9
              "01010" when "11001", -- t[25] = 10
              "01011" when "11010", -- t[26] = 11
              "01100" when "11011", -- t[27] = 12
              "01100" when "11100", -- t[28] = 12
              "01101" when "11101", -- t[29] = 13
              "01110" when "11110", -- t[30] = 14
              "01111" when "11111", -- t[31] = 15
              "-----" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_9 is
  port ( nY2    : in  std_logic_vector(3 downto 0);
         nExpY2 : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_9 is
begin

  with nY2 select
    nExpY2 <= "0000" when "0000", -- t[0] = 0
              "0000" when "0001", -- t[1] = 0
              "0000" when "0010", -- t[2] = 0
              "0000" when "0011", -- t[3] = 0
              "0001" when "0100", -- t[4] = 1
              "0001" when "0101", -- t[5] = 1
              "0001" when "0110", -- t[6] = 1
              "0010" when "0111", -- t[7] = 2
              "0010" when "1000", -- t[8] = 2
              "0011" when "1001", -- t[9] = 3
              "0011" when "1010", -- t[10] = 3
              "0100" when "1011", -- t[11] = 4
              "0101" when "1100", -- t[12] = 5
              "0101" when "1101", -- t[13] = 5
              "0110" when "1110", -- t[14] = 6
              "0111" when "1111", -- t[15] = 7
              "----" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_10 is
  port ( nY2    : in  std_logic_vector(4 downto 0);
         nExpY2 : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_10 is
begin

  with nY2 select
    nExpY2 <= "00000" when "00000", -- t[0] = 0
              "00000" when "00001", -- t[1] = 0
              "00000" when "00010", -- t[2] = 0
              "00000" when "00011", -- t[3] = 0
              "00000" when "00100", -- t[4] = 0
              "00000" when "00101", -- t[5] = 0
              "00001" when "00110", -- t[6] = 1
              "00001" when "00111", -- t[7] = 1
              "00001" when "01000", -- t[8] = 1
              "00001" when "01001", -- t[9] = 1
              "00010" when "01010", -- t[10] = 2
              "00010" when "01011", -- t[11] = 2
              "00010" when "01100", -- t[12] = 2
              "00011" when "01101", -- t[13] = 3
              "00011" when "01110", -- t[14] = 3
              "00100" when "01111", -- t[15] = 4
              "00100" when "10000", -- t[16] = 4
              "00101" when "10001", -- t[17] = 5
              "00101" when "10010", -- t[18] = 5
              "00110" when "10011", -- t[19] = 6
              "00110" when "10100", -- t[20] = 6
              "00111" when "10101", -- t[21] = 7
              "01000" when "10110", -- t[22] = 8
              "01000" when "10111", -- t[23] = 8
              "01001" when "11000", -- t[24] = 9
              "01010" when "11001", -- t[25] = 10
              "01011" when "11010", -- t[26] = 11
              "01011" when "11011", -- t[27] = 11
              "01100" when "11100", -- t[28] = 12
              "01101" when "11101", -- t[29] = 13
              "01110" when "11110", -- t[30] = 14
              "01111" when "11111", -- t[31] = 15
              "-----" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_11 is
  port ( nY2    : in  std_logic_vector(5 downto 0);
         nExpY2 : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_11 is
begin

  with nY2 select
    nExpY2 <= "000000" when "000000", -- t[0] = 0
              "000000" when "000001", -- t[1] = 0
              "000000" when "000010", -- t[2] = 0
              "000000" when "000011", -- t[3] = 0
              "000000" when "000100", -- t[4] = 0
              "000000" when "000101", -- t[5] = 0
              "000000" when "000110", -- t[6] = 0
              "000000" when "000111", -- t[7] = 0
              "000001" when "001000", -- t[8] = 1
              "000001" when "001001", -- t[9] = 1
              "000001" when "001010", -- t[10] = 1
              "000001" when "001011", -- t[11] = 1
              "000001" when "001100", -- t[12] = 1
              "000001" when "001101", -- t[13] = 1
              "000010" when "001110", -- t[14] = 2
              "000010" when "001111", -- t[15] = 2
              "000010" when "010000", -- t[16] = 2
              "000010" when "010001", -- t[17] = 2
              "000011" when "010010", -- t[18] = 3
              "000011" when "010011", -- t[19] = 3
              "000011" when "010100", -- t[20] = 3
              "000011" when "010101", -- t[21] = 3
              "000100" when "010110", -- t[22] = 4
              "000100" when "010111", -- t[23] = 4
              "000101" when "011000", -- t[24] = 5
              "000101" when "011001", -- t[25] = 5
              "000101" when "011010", -- t[26] = 5
              "000110" when "011011", -- t[27] = 6
              "000110" when "011100", -- t[28] = 6
              "000111" when "011101", -- t[29] = 7
              "000111" when "011110", -- t[30] = 7
              "001000" when "011111", -- t[31] = 8
              "001000" when "100000", -- t[32] = 8
              "001001" when "100001", -- t[33] = 9
              "001001" when "100010", -- t[34] = 9
              "001010" when "100011", -- t[35] = 10
              "001010" when "100100", -- t[36] = 10
              "001011" when "100101", -- t[37] = 11
              "001011" when "100110", -- t[38] = 11
              "001100" when "100111", -- t[39] = 12
              "001101" when "101000", -- t[40] = 13
              "001101" when "101001", -- t[41] = 13
              "001110" when "101010", -- t[42] = 14
              "001111" when "101011", -- t[43] = 15
              "001111" when "101100", -- t[44] = 15
              "010000" when "101101", -- t[45] = 16
              "010001" when "101110", -- t[46] = 17
              "010001" when "101111", -- t[47] = 17
              "010010" when "110000", -- t[48] = 18
              "010011" when "110001", -- t[49] = 19
              "010100" when "110010", -- t[50] = 20
              "010100" when "110011", -- t[51] = 20
              "010101" when "110100", -- t[52] = 21
              "010110" when "110101", -- t[53] = 22
              "010111" when "110110", -- t[54] = 23
              "011000" when "110111", -- t[55] = 24
              "011001" when "111000", -- t[56] = 25
              "011010" when "111001", -- t[57] = 26
              "011011" when "111010", -- t[58] = 27
              "011011" when "111011", -- t[59] = 27
              "011100" when "111100", -- t[60] = 28
              "011101" when "111101", -- t[61] = 29
              "011110" when "111110", -- t[62] = 30
              "011111" when "111111", -- t[63] = 31
              "------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_12 is
  port ( nY2    : in  std_logic_vector(4 downto 0);
         nExpY2 : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_12 is
begin

  with nY2 select
    nExpY2 <= "00000" when "00000", -- t[0] = 0
              "00000" when "00001", -- t[1] = 0
              "00000" when "00010", -- t[2] = 0
              "00000" when "00011", -- t[3] = 0
              "00000" when "00100", -- t[4] = 0
              "00000" when "00101", -- t[5] = 0
              "00001" when "00110", -- t[6] = 1
              "00001" when "00111", -- t[7] = 1
              "00001" when "01000", -- t[8] = 1
              "00001" when "01001", -- t[9] = 1
              "00010" when "01010", -- t[10] = 2
              "00010" when "01011", -- t[11] = 2
              "00010" when "01100", -- t[12] = 2
              "00011" when "01101", -- t[13] = 3
              "00011" when "01110", -- t[14] = 3
              "00100" when "01111", -- t[15] = 4
              "00100" when "10000", -- t[16] = 4
              "00101" when "10001", -- t[17] = 5
              "00101" when "10010", -- t[18] = 5
              "00110" when "10011", -- t[19] = 6
              "00110" when "10100", -- t[20] = 6
              "00111" when "10101", -- t[21] = 7
              "01000" when "10110", -- t[22] = 8
              "01000" when "10111", -- t[23] = 8
              "01001" when "11000", -- t[24] = 9
              "01010" when "11001", -- t[25] = 10
              "01011" when "11010", -- t[26] = 11
              "01011" when "11011", -- t[27] = 11
              "01100" when "11100", -- t[28] = 12
              "01101" when "11101", -- t[29] = 13
              "01110" when "11110", -- t[30] = 14
              "01111" when "11111", -- t[31] = 15
              "-----" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_13 is
  port ( nY2    : in  std_logic_vector(5 downto 0);
         nExpY2 : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_13 is
begin

  with nY2 select
    nExpY2 <= "000000" when "000000", -- t[0] = 0
              "000000" when "000001", -- t[1] = 0
              "000000" when "000010", -- t[2] = 0
              "000000" when "000011", -- t[3] = 0
              "000000" when "000100", -- t[4] = 0
              "000000" when "000101", -- t[5] = 0
              "000000" when "000110", -- t[6] = 0
              "000000" when "000111", -- t[7] = 0
              "000001" when "001000", -- t[8] = 1
              "000001" when "001001", -- t[9] = 1
              "000001" when "001010", -- t[10] = 1
              "000001" when "001011", -- t[11] = 1
              "000001" when "001100", -- t[12] = 1
              "000001" when "001101", -- t[13] = 1
              "000010" when "001110", -- t[14] = 2
              "000010" when "001111", -- t[15] = 2
              "000010" when "010000", -- t[16] = 2
              "000010" when "010001", -- t[17] = 2
              "000011" when "010010", -- t[18] = 3
              "000011" when "010011", -- t[19] = 3
              "000011" when "010100", -- t[20] = 3
              "000011" when "010101", -- t[21] = 3
              "000100" when "010110", -- t[22] = 4
              "000100" when "010111", -- t[23] = 4
              "000101" when "011000", -- t[24] = 5
              "000101" when "011001", -- t[25] = 5
              "000101" when "011010", -- t[26] = 5
              "000110" when "011011", -- t[27] = 6
              "000110" when "011100", -- t[28] = 6
              "000111" when "011101", -- t[29] = 7
              "000111" when "011110", -- t[30] = 7
              "001000" when "011111", -- t[31] = 8
              "001000" when "100000", -- t[32] = 8
              "001001" when "100001", -- t[33] = 9
              "001001" when "100010", -- t[34] = 9
              "001010" when "100011", -- t[35] = 10
              "001010" when "100100", -- t[36] = 10
              "001011" when "100101", -- t[37] = 11
              "001011" when "100110", -- t[38] = 11
              "001100" when "100111", -- t[39] = 12
              "001101" when "101000", -- t[40] = 13
              "001101" when "101001", -- t[41] = 13
              "001110" when "101010", -- t[42] = 14
              "001110" when "101011", -- t[43] = 14
              "001111" when "101100", -- t[44] = 15
              "010000" when "101101", -- t[45] = 16
              "010001" when "101110", -- t[46] = 17
              "010001" when "101111", -- t[47] = 17
              "010010" when "110000", -- t[48] = 18
              "010011" when "110001", -- t[49] = 19
              "010100" when "110010", -- t[50] = 20
              "010100" when "110011", -- t[51] = 20
              "010101" when "110100", -- t[52] = 21
              "010110" when "110101", -- t[53] = 22
              "010111" when "110110", -- t[54] = 23
              "011000" when "110111", -- t[55] = 24
              "011001" when "111000", -- t[56] = 25
              "011010" when "111001", -- t[57] = 26
              "011010" when "111010", -- t[58] = 26
              "011011" when "111011", -- t[59] = 27
              "011100" when "111100", -- t[60] = 28
              "011101" when "111101", -- t[61] = 29
              "011110" when "111110", -- t[62] = 30
              "011111" when "111111", -- t[63] = 31
              "------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_14 is
  port ( nY2    : in  std_logic_vector(6 downto 0);
         nExpY2 : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_14 is
begin

  with nY2 select
    nExpY2 <= "0000000" when "0000000", -- t[0] = 0
              "0000000" when "0000001", -- t[1] = 0
              "0000000" when "0000010", -- t[2] = 0
              "0000000" when "0000011", -- t[3] = 0
              "0000000" when "0000100", -- t[4] = 0
              "0000000" when "0000101", -- t[5] = 0
              "0000000" when "0000110", -- t[6] = 0
              "0000000" when "0000111", -- t[7] = 0
              "0000000" when "0001000", -- t[8] = 0
              "0000000" when "0001001", -- t[9] = 0
              "0000000" when "0001010", -- t[10] = 0
              "0000000" when "0001011", -- t[11] = 0
              "0000001" when "0001100", -- t[12] = 1
              "0000001" when "0001101", -- t[13] = 1
              "0000001" when "0001110", -- t[14] = 1
              "0000001" when "0001111", -- t[15] = 1
              "0000001" when "0010000", -- t[16] = 1
              "0000001" when "0010001", -- t[17] = 1
              "0000001" when "0010010", -- t[18] = 1
              "0000001" when "0010011", -- t[19] = 1
              "0000010" when "0010100", -- t[20] = 2
              "0000010" when "0010101", -- t[21] = 2
              "0000010" when "0010110", -- t[22] = 2
              "0000010" when "0010111", -- t[23] = 2
              "0000010" when "0011000", -- t[24] = 2
              "0000010" when "0011001", -- t[25] = 2
              "0000011" when "0011010", -- t[26] = 3
              "0000011" when "0011011", -- t[27] = 3
              "0000011" when "0011100", -- t[28] = 3
              "0000011" when "0011101", -- t[29] = 3
              "0000100" when "0011110", -- t[30] = 4
              "0000100" when "0011111", -- t[31] = 4
              "0000100" when "0100000", -- t[32] = 4
              "0000100" when "0100001", -- t[33] = 4
              "0000101" when "0100010", -- t[34] = 5
              "0000101" when "0100011", -- t[35] = 5
              "0000101" when "0100100", -- t[36] = 5
              "0000101" when "0100101", -- t[37] = 5
              "0000110" when "0100110", -- t[38] = 6
              "0000110" when "0100111", -- t[39] = 6
              "0000110" when "0101000", -- t[40] = 6
              "0000111" when "0101001", -- t[41] = 7
              "0000111" when "0101010", -- t[42] = 7
              "0000111" when "0101011", -- t[43] = 7
              "0001000" when "0101100", -- t[44] = 8
              "0001000" when "0101101", -- t[45] = 8
              "0001000" when "0101110", -- t[46] = 8
              "0001001" when "0101111", -- t[47] = 9
              "0001001" when "0110000", -- t[48] = 9
              "0001001" when "0110001", -- t[49] = 9
              "0001010" when "0110010", -- t[50] = 10
              "0001010" when "0110011", -- t[51] = 10
              "0001011" when "0110100", -- t[52] = 11
              "0001011" when "0110101", -- t[53] = 11
              "0001011" when "0110110", -- t[54] = 11
              "0001100" when "0110111", -- t[55] = 12
              "0001100" when "0111000", -- t[56] = 12
              "0001101" when "0111001", -- t[57] = 13
              "0001101" when "0111010", -- t[58] = 13
              "0001110" when "0111011", -- t[59] = 14
              "0001110" when "0111100", -- t[60] = 14
              "0001111" when "0111101", -- t[61] = 15
              "0001111" when "0111110", -- t[62] = 15
              "0010000" when "0111111", -- t[63] = 16
              "0010000" when "1000000", -- t[64] = 16
              "0010001" when "1000001", -- t[65] = 17
              "0010001" when "1000010", -- t[66] = 17
              "0010010" when "1000011", -- t[67] = 18
              "0010010" when "1000100", -- t[68] = 18
              "0010011" when "1000101", -- t[69] = 19
              "0010011" when "1000110", -- t[70] = 19
              "0010100" when "1000111", -- t[71] = 20
              "0010100" when "1001000", -- t[72] = 20
              "0010101" when "1001001", -- t[73] = 21
              "0010101" when "1001010", -- t[74] = 21
              "0010110" when "1001011", -- t[75] = 22
              "0010111" when "1001100", -- t[76] = 23
              "0010111" when "1001101", -- t[77] = 23
              "0011000" when "1001110", -- t[78] = 24
              "0011000" when "1001111", -- t[79] = 24
              "0011001" when "1010000", -- t[80] = 25
              "0011010" when "1010001", -- t[81] = 26
              "0011010" when "1010010", -- t[82] = 26
              "0011011" when "1010011", -- t[83] = 27
              "0011100" when "1010100", -- t[84] = 28
              "0011100" when "1010101", -- t[85] = 28
              "0011101" when "1010110", -- t[86] = 29
              "0011110" when "1010111", -- t[87] = 30
              "0011110" when "1011000", -- t[88] = 30
              "0011111" when "1011001", -- t[89] = 31
              "0100000" when "1011010", -- t[90] = 32
              "0100000" when "1011011", -- t[91] = 32
              "0100001" when "1011100", -- t[92] = 33
              "0100010" when "1011101", -- t[93] = 34
              "0100011" when "1011110", -- t[94] = 35
              "0100011" when "1011111", -- t[95] = 35
              "0100100" when "1100000", -- t[96] = 36
              "0100101" when "1100001", -- t[97] = 37
              "0100110" when "1100010", -- t[98] = 38
              "0100110" when "1100011", -- t[99] = 38
              "0100111" when "1100100", -- t[100] = 39
              "0101000" when "1100101", -- t[101] = 40
              "0101001" when "1100110", -- t[102] = 41
              "0101010" when "1100111", -- t[103] = 42
              "0101010" when "1101000", -- t[104] = 42
              "0101011" when "1101001", -- t[105] = 43
              "0101100" when "1101010", -- t[106] = 44
              "0101101" when "1101011", -- t[107] = 45
              "0101110" when "1101100", -- t[108] = 46
              "0101111" when "1101101", -- t[109] = 47
              "0101111" when "1101110", -- t[110] = 47
              "0110000" when "1101111", -- t[111] = 48
              "0110001" when "1110000", -- t[112] = 49
              "0110010" when "1110001", -- t[113] = 50
              "0110011" when "1110010", -- t[114] = 51
              "0110100" when "1110011", -- t[115] = 52
              "0110101" when "1110100", -- t[116] = 53
              "0110110" when "1110101", -- t[117] = 54
              "0110111" when "1110110", -- t[118] = 55
              "0111000" when "1110111", -- t[119] = 56
              "0111001" when "1111000", -- t[120] = 57
              "0111001" when "1111001", -- t[121] = 57
              "0111010" when "1111010", -- t[122] = 58
              "0111011" when "1111011", -- t[123] = 59
              "0111100" when "1111100", -- t[124] = 60
              "0111101" when "1111101", -- t[125] = 61
              "0111110" when "1111110", -- t[126] = 62
              "0111111" when "1111111", -- t[127] = 63
              "-------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_15 is
  port ( nY2    : in  std_logic_vector(5 downto 0);
         nExpY2 : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_15 is
begin

  with nY2 select
    nExpY2 <= "000000" when "000000", -- t[0] = 0
              "000000" when "000001", -- t[1] = 0
              "000000" when "000010", -- t[2] = 0
              "000000" when "000011", -- t[3] = 0
              "000000" when "000100", -- t[4] = 0
              "000000" when "000101", -- t[5] = 0
              "000000" when "000110", -- t[6] = 0
              "000000" when "000111", -- t[7] = 0
              "000001" when "001000", -- t[8] = 1
              "000001" when "001001", -- t[9] = 1
              "000001" when "001010", -- t[10] = 1
              "000001" when "001011", -- t[11] = 1
              "000001" when "001100", -- t[12] = 1
              "000001" when "001101", -- t[13] = 1
              "000010" when "001110", -- t[14] = 2
              "000010" when "001111", -- t[15] = 2
              "000010" when "010000", -- t[16] = 2
              "000010" when "010001", -- t[17] = 2
              "000011" when "010010", -- t[18] = 3
              "000011" when "010011", -- t[19] = 3
              "000011" when "010100", -- t[20] = 3
              "000011" when "010101", -- t[21] = 3
              "000100" when "010110", -- t[22] = 4
              "000100" when "010111", -- t[23] = 4
              "000101" when "011000", -- t[24] = 5
              "000101" when "011001", -- t[25] = 5
              "000101" when "011010", -- t[26] = 5
              "000110" when "011011", -- t[27] = 6
              "000110" when "011100", -- t[28] = 6
              "000111" when "011101", -- t[29] = 7
              "000111" when "011110", -- t[30] = 7
              "001000" when "011111", -- t[31] = 8
              "001000" when "100000", -- t[32] = 8
              "001001" when "100001", -- t[33] = 9
              "001001" when "100010", -- t[34] = 9
              "001010" when "100011", -- t[35] = 10
              "001010" when "100100", -- t[36] = 10
              "001011" when "100101", -- t[37] = 11
              "001011" when "100110", -- t[38] = 11
              "001100" when "100111", -- t[39] = 12
              "001101" when "101000", -- t[40] = 13
              "001101" when "101001", -- t[41] = 13
              "001110" when "101010", -- t[42] = 14
              "001110" when "101011", -- t[43] = 14
              "001111" when "101100", -- t[44] = 15
              "010000" when "101101", -- t[45] = 16
              "010001" when "101110", -- t[46] = 17
              "010001" when "101111", -- t[47] = 17
              "010010" when "110000", -- t[48] = 18
              "010011" when "110001", -- t[49] = 19
              "010100" when "110010", -- t[50] = 20
              "010100" when "110011", -- t[51] = 20
              "010101" when "110100", -- t[52] = 21
              "010110" when "110101", -- t[53] = 22
              "010111" when "110110", -- t[54] = 23
              "011000" when "110111", -- t[55] = 24
              "011001" when "111000", -- t[56] = 25
              "011001" when "111001", -- t[57] = 25
              "011010" when "111010", -- t[58] = 26
              "011011" when "111011", -- t[59] = 27
              "011100" when "111100", -- t[60] = 28
              "011101" when "111101", -- t[61] = 29
              "011110" when "111110", -- t[62] = 30
              "011111" when "111111", -- t[63] = 31
              "------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_16 is
  port ( nY2    : in  std_logic_vector(6 downto 0);
         nExpY2 : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_16 is
begin

  with nY2 select
    nExpY2 <= "0000000" when "0000000", -- t[0] = 0
              "0000000" when "0000001", -- t[1] = 0
              "0000000" when "0000010", -- t[2] = 0
              "0000000" when "0000011", -- t[3] = 0
              "0000000" when "0000100", -- t[4] = 0
              "0000000" when "0000101", -- t[5] = 0
              "0000000" when "0000110", -- t[6] = 0
              "0000000" when "0000111", -- t[7] = 0
              "0000000" when "0001000", -- t[8] = 0
              "0000000" when "0001001", -- t[9] = 0
              "0000000" when "0001010", -- t[10] = 0
              "0000000" when "0001011", -- t[11] = 0
              "0000001" when "0001100", -- t[12] = 1
              "0000001" when "0001101", -- t[13] = 1
              "0000001" when "0001110", -- t[14] = 1
              "0000001" when "0001111", -- t[15] = 1
              "0000001" when "0010000", -- t[16] = 1
              "0000001" when "0010001", -- t[17] = 1
              "0000001" when "0010010", -- t[18] = 1
              "0000001" when "0010011", -- t[19] = 1
              "0000010" when "0010100", -- t[20] = 2
              "0000010" when "0010101", -- t[21] = 2
              "0000010" when "0010110", -- t[22] = 2
              "0000010" when "0010111", -- t[23] = 2
              "0000010" when "0011000", -- t[24] = 2
              "0000010" when "0011001", -- t[25] = 2
              "0000011" when "0011010", -- t[26] = 3
              "0000011" when "0011011", -- t[27] = 3
              "0000011" when "0011100", -- t[28] = 3
              "0000011" when "0011101", -- t[29] = 3
              "0000100" when "0011110", -- t[30] = 4
              "0000100" when "0011111", -- t[31] = 4
              "0000100" when "0100000", -- t[32] = 4
              "0000100" when "0100001", -- t[33] = 4
              "0000101" when "0100010", -- t[34] = 5
              "0000101" when "0100011", -- t[35] = 5
              "0000101" when "0100100", -- t[36] = 5
              "0000101" when "0100101", -- t[37] = 5
              "0000110" when "0100110", -- t[38] = 6
              "0000110" when "0100111", -- t[39] = 6
              "0000110" when "0101000", -- t[40] = 6
              "0000111" when "0101001", -- t[41] = 7
              "0000111" when "0101010", -- t[42] = 7
              "0000111" when "0101011", -- t[43] = 7
              "0001000" when "0101100", -- t[44] = 8
              "0001000" when "0101101", -- t[45] = 8
              "0001000" when "0101110", -- t[46] = 8
              "0001001" when "0101111", -- t[47] = 9
              "0001001" when "0110000", -- t[48] = 9
              "0001001" when "0110001", -- t[49] = 9
              "0001010" when "0110010", -- t[50] = 10
              "0001010" when "0110011", -- t[51] = 10
              "0001011" when "0110100", -- t[52] = 11
              "0001011" when "0110101", -- t[53] = 11
              "0001011" when "0110110", -- t[54] = 11
              "0001100" when "0110111", -- t[55] = 12
              "0001100" when "0111000", -- t[56] = 12
              "0001101" when "0111001", -- t[57] = 13
              "0001101" when "0111010", -- t[58] = 13
              "0001110" when "0111011", -- t[59] = 14
              "0001110" when "0111100", -- t[60] = 14
              "0001111" when "0111101", -- t[61] = 15
              "0001111" when "0111110", -- t[62] = 15
              "0010000" when "0111111", -- t[63] = 16
              "0010000" when "1000000", -- t[64] = 16
              "0010001" when "1000001", -- t[65] = 17
              "0010001" when "1000010", -- t[66] = 17
              "0010010" when "1000011", -- t[67] = 18
              "0010010" when "1000100", -- t[68] = 18
              "0010011" when "1000101", -- t[69] = 19
              "0010011" when "1000110", -- t[70] = 19
              "0010100" when "1000111", -- t[71] = 20
              "0010100" when "1001000", -- t[72] = 20
              "0010101" when "1001001", -- t[73] = 21
              "0010101" when "1001010", -- t[74] = 21
              "0010110" when "1001011", -- t[75] = 22
              "0010111" when "1001100", -- t[76] = 23
              "0010111" when "1001101", -- t[77] = 23
              "0011000" when "1001110", -- t[78] = 24
              "0011000" when "1001111", -- t[79] = 24
              "0011001" when "1010000", -- t[80] = 25
              "0011010" when "1010001", -- t[81] = 26
              "0011010" when "1010010", -- t[82] = 26
              "0011011" when "1010011", -- t[83] = 27
              "0011100" when "1010100", -- t[84] = 28
              "0011100" when "1010101", -- t[85] = 28
              "0011101" when "1010110", -- t[86] = 29
              "0011110" when "1010111", -- t[87] = 30
              "0011110" when "1011000", -- t[88] = 30
              "0011111" when "1011001", -- t[89] = 31
              "0100000" when "1011010", -- t[90] = 32
              "0100000" when "1011011", -- t[91] = 32
              "0100001" when "1011100", -- t[92] = 33
              "0100010" when "1011101", -- t[93] = 34
              "0100011" when "1011110", -- t[94] = 35
              "0100011" when "1011111", -- t[95] = 35
              "0100100" when "1100000", -- t[96] = 36
              "0100101" when "1100001", -- t[97] = 37
              "0100110" when "1100010", -- t[98] = 38
              "0100110" when "1100011", -- t[99] = 38
              "0100111" when "1100100", -- t[100] = 39
              "0101000" when "1100101", -- t[101] = 40
              "0101001" when "1100110", -- t[102] = 41
              "0101010" when "1100111", -- t[103] = 42
              "0101010" when "1101000", -- t[104] = 42
              "0101011" when "1101001", -- t[105] = 43
              "0101100" when "1101010", -- t[106] = 44
              "0101101" when "1101011", -- t[107] = 45
              "0101110" when "1101100", -- t[108] = 46
              "0101111" when "1101101", -- t[109] = 47
              "0101111" when "1101110", -- t[110] = 47
              "0110000" when "1101111", -- t[111] = 48
              "0110001" when "1110000", -- t[112] = 49
              "0110010" when "1110001", -- t[113] = 50
              "0110011" when "1110010", -- t[114] = 51
              "0110100" when "1110011", -- t[115] = 52
              "0110101" when "1110100", -- t[116] = 53
              "0110110" when "1110101", -- t[117] = 54
              "0110111" when "1110110", -- t[118] = 55
              "0110111" when "1110111", -- t[119] = 55
              "0111000" when "1111000", -- t[120] = 56
              "0111001" when "1111001", -- t[121] = 57
              "0111010" when "1111010", -- t[122] = 58
              "0111011" when "1111011", -- t[123] = 59
              "0111100" when "1111100", -- t[124] = 60
              "0111101" when "1111101", -- t[125] = 61
              "0111110" when "1111110", -- t[126] = 62
              "0111111" when "1111111", -- t[127] = 63
              "-------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_17 is
  port ( nY2    : in  std_logic_vector(7 downto 0);
         nExpY2 : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_17 is
begin

  with nY2 select
    nExpY2 <= "00000000" when "00000000", -- t[0] = 0
              "00000000" when "00000001", -- t[1] = 0
              "00000000" when "00000010", -- t[2] = 0
              "00000000" when "00000011", -- t[3] = 0
              "00000000" when "00000100", -- t[4] = 0
              "00000000" when "00000101", -- t[5] = 0
              "00000000" when "00000110", -- t[6] = 0
              "00000000" when "00000111", -- t[7] = 0
              "00000000" when "00001000", -- t[8] = 0
              "00000000" when "00001001", -- t[9] = 0
              "00000000" when "00001010", -- t[10] = 0
              "00000000" when "00001011", -- t[11] = 0
              "00000000" when "00001100", -- t[12] = 0
              "00000000" when "00001101", -- t[13] = 0
              "00000000" when "00001110", -- t[14] = 0
              "00000000" when "00001111", -- t[15] = 0
              "00000001" when "00010000", -- t[16] = 1
              "00000001" when "00010001", -- t[17] = 1
              "00000001" when "00010010", -- t[18] = 1
              "00000001" when "00010011", -- t[19] = 1
              "00000001" when "00010100", -- t[20] = 1
              "00000001" when "00010101", -- t[21] = 1
              "00000001" when "00010110", -- t[22] = 1
              "00000001" when "00010111", -- t[23] = 1
              "00000001" when "00011000", -- t[24] = 1
              "00000001" when "00011001", -- t[25] = 1
              "00000001" when "00011010", -- t[26] = 1
              "00000001" when "00011011", -- t[27] = 1
              "00000010" when "00011100", -- t[28] = 2
              "00000010" when "00011101", -- t[29] = 2
              "00000010" when "00011110", -- t[30] = 2
              "00000010" when "00011111", -- t[31] = 2
              "00000010" when "00100000", -- t[32] = 2
              "00000010" when "00100001", -- t[33] = 2
              "00000010" when "00100010", -- t[34] = 2
              "00000010" when "00100011", -- t[35] = 2
              "00000011" when "00100100", -- t[36] = 3
              "00000011" when "00100101", -- t[37] = 3
              "00000011" when "00100110", -- t[38] = 3
              "00000011" when "00100111", -- t[39] = 3
              "00000011" when "00101000", -- t[40] = 3
              "00000011" when "00101001", -- t[41] = 3
              "00000011" when "00101010", -- t[42] = 3
              "00000100" when "00101011", -- t[43] = 4
              "00000100" when "00101100", -- t[44] = 4
              "00000100" when "00101101", -- t[45] = 4
              "00000100" when "00101110", -- t[46] = 4
              "00000100" when "00101111", -- t[47] = 4
              "00000101" when "00110000", -- t[48] = 5
              "00000101" when "00110001", -- t[49] = 5
              "00000101" when "00110010", -- t[50] = 5
              "00000101" when "00110011", -- t[51] = 5
              "00000101" when "00110100", -- t[52] = 5
              "00000101" when "00110101", -- t[53] = 5
              "00000110" when "00110110", -- t[54] = 6
              "00000110" when "00110111", -- t[55] = 6
              "00000110" when "00111000", -- t[56] = 6
              "00000110" when "00111001", -- t[57] = 6
              "00000111" when "00111010", -- t[58] = 7
              "00000111" when "00111011", -- t[59] = 7
              "00000111" when "00111100", -- t[60] = 7
              "00000111" when "00111101", -- t[61] = 7
              "00001000" when "00111110", -- t[62] = 8
              "00001000" when "00111111", -- t[63] = 8
              "00001000" when "01000000", -- t[64] = 8
              "00001000" when "01000001", -- t[65] = 8
              "00001001" when "01000010", -- t[66] = 9
              "00001001" when "01000011", -- t[67] = 9
              "00001001" when "01000100", -- t[68] = 9
              "00001001" when "01000101", -- t[69] = 9
              "00001010" when "01000110", -- t[70] = 10
              "00001010" when "01000111", -- t[71] = 10
              "00001010" when "01001000", -- t[72] = 10
              "00001010" when "01001001", -- t[73] = 10
              "00001011" when "01001010", -- t[74] = 11
              "00001011" when "01001011", -- t[75] = 11
              "00001011" when "01001100", -- t[76] = 11
              "00001100" when "01001101", -- t[77] = 12
              "00001100" when "01001110", -- t[78] = 12
              "00001100" when "01001111", -- t[79] = 12
              "00001101" when "01010000", -- t[80] = 13
              "00001101" when "01010001", -- t[81] = 13
              "00001101" when "01010010", -- t[82] = 13
              "00001101" when "01010011", -- t[83] = 13
              "00001110" when "01010100", -- t[84] = 14
              "00001110" when "01010101", -- t[85] = 14
              "00001110" when "01010110", -- t[86] = 14
              "00001111" when "01010111", -- t[87] = 15
              "00001111" when "01011000", -- t[88] = 15
              "00001111" when "01011001", -- t[89] = 15
              "00010000" when "01011010", -- t[90] = 16
              "00010000" when "01011011", -- t[91] = 16
              "00010001" when "01011100", -- t[92] = 17
              "00010001" when "01011101", -- t[93] = 17
              "00010001" when "01011110", -- t[94] = 17
              "00010010" when "01011111", -- t[95] = 18
              "00010010" when "01100000", -- t[96] = 18
              "00010010" when "01100001", -- t[97] = 18
              "00010011" when "01100010", -- t[98] = 19
              "00010011" when "01100011", -- t[99] = 19
              "00010100" when "01100100", -- t[100] = 20
              "00010100" when "01100101", -- t[101] = 20
              "00010100" when "01100110", -- t[102] = 20
              "00010101" when "01100111", -- t[103] = 21
              "00010101" when "01101000", -- t[104] = 21
              "00010110" when "01101001", -- t[105] = 22
              "00010110" when "01101010", -- t[106] = 22
              "00010110" when "01101011", -- t[107] = 22
              "00010111" when "01101100", -- t[108] = 23
              "00010111" when "01101101", -- t[109] = 23
              "00011000" when "01101110", -- t[110] = 24
              "00011000" when "01101111", -- t[111] = 24
              "00011001" when "01110000", -- t[112] = 25
              "00011001" when "01110001", -- t[113] = 25
              "00011001" when "01110010", -- t[114] = 25
              "00011010" when "01110011", -- t[115] = 26
              "00011010" when "01110100", -- t[116] = 26
              "00011011" when "01110101", -- t[117] = 27
              "00011011" when "01110110", -- t[118] = 27
              "00011100" when "01110111", -- t[119] = 28
              "00011100" when "01111000", -- t[120] = 28
              "00011101" when "01111001", -- t[121] = 29
              "00011101" when "01111010", -- t[122] = 29
              "00011110" when "01111011", -- t[123] = 30
              "00011110" when "01111100", -- t[124] = 30
              "00011111" when "01111101", -- t[125] = 31
              "00011111" when "01111110", -- t[126] = 31
              "00100000" when "01111111", -- t[127] = 32
              "00100000" when "10000000", -- t[128] = 32
              "00100001" when "10000001", -- t[129] = 33
              "00100001" when "10000010", -- t[130] = 33
              "00100010" when "10000011", -- t[131] = 34
              "00100010" when "10000100", -- t[132] = 34
              "00100011" when "10000101", -- t[133] = 35
              "00100011" when "10000110", -- t[134] = 35
              "00100100" when "10000111", -- t[135] = 36
              "00100100" when "10001000", -- t[136] = 36
              "00100101" when "10001001", -- t[137] = 37
              "00100101" when "10001010", -- t[138] = 37
              "00100110" when "10001011", -- t[139] = 38
              "00100110" when "10001100", -- t[140] = 38
              "00100111" when "10001101", -- t[141] = 39
              "00100111" when "10001110", -- t[142] = 39
              "00101000" when "10001111", -- t[143] = 40
              "00101001" when "10010000", -- t[144] = 41
              "00101001" when "10010001", -- t[145] = 41
              "00101010" when "10010010", -- t[146] = 42
              "00101010" when "10010011", -- t[147] = 42
              "00101011" when "10010100", -- t[148] = 43
              "00101011" when "10010101", -- t[149] = 43
              "00101100" when "10010110", -- t[150] = 44
              "00101101" when "10010111", -- t[151] = 45
              "00101101" when "10011000", -- t[152] = 45
              "00101110" when "10011001", -- t[153] = 46
              "00101110" when "10011010", -- t[154] = 46
              "00101111" when "10011011", -- t[155] = 47
              "00110000" when "10011100", -- t[156] = 48
              "00110000" when "10011101", -- t[157] = 48
              "00110001" when "10011110", -- t[158] = 49
              "00110001" when "10011111", -- t[159] = 49
              "00110010" when "10100000", -- t[160] = 50
              "00110011" when "10100001", -- t[161] = 51
              "00110011" when "10100010", -- t[162] = 51
              "00110100" when "10100011", -- t[163] = 52
              "00110101" when "10100100", -- t[164] = 53
              "00110101" when "10100101", -- t[165] = 53
              "00110110" when "10100110", -- t[166] = 54
              "00110111" when "10100111", -- t[167] = 55
              "00110111" when "10101000", -- t[168] = 55
              "00111000" when "10101001", -- t[169] = 56
              "00111001" when "10101010", -- t[170] = 57
              "00111001" when "10101011", -- t[171] = 57
              "00111010" when "10101100", -- t[172] = 58
              "00111011" when "10101101", -- t[173] = 59
              "00111011" when "10101110", -- t[174] = 59
              "00111100" when "10101111", -- t[175] = 60
              "00111101" when "10110000", -- t[176] = 61
              "00111101" when "10110001", -- t[177] = 61
              "00111110" when "10110010", -- t[178] = 62
              "00111111" when "10110011", -- t[179] = 63
              "00111111" when "10110100", -- t[180] = 63
              "01000000" when "10110101", -- t[181] = 64
              "01000001" when "10110110", -- t[182] = 65
              "01000010" when "10110111", -- t[183] = 66
              "01000010" when "10111000", -- t[184] = 66
              "01000011" when "10111001", -- t[185] = 67
              "01000100" when "10111010", -- t[186] = 68
              "01000100" when "10111011", -- t[187] = 68
              "01000101" when "10111100", -- t[188] = 69
              "01000110" when "10111101", -- t[189] = 70
              "01000111" when "10111110", -- t[190] = 71
              "01000111" when "10111111", -- t[191] = 71
              "01001000" when "11000000", -- t[192] = 72
              "01001001" when "11000001", -- t[193] = 73
              "01001010" when "11000010", -- t[194] = 74
              "01001010" when "11000011", -- t[195] = 74
              "01001011" when "11000100", -- t[196] = 75
              "01001100" when "11000101", -- t[197] = 76
              "01001101" when "11000110", -- t[198] = 77
              "01001110" when "11000111", -- t[199] = 78
              "01001110" when "11001000", -- t[200] = 78
              "01001111" when "11001001", -- t[201] = 79
              "01010000" when "11001010", -- t[202] = 80
              "01010001" when "11001011", -- t[203] = 81
              "01010001" when "11001100", -- t[204] = 81
              "01010010" when "11001101", -- t[205] = 82
              "01010011" when "11001110", -- t[206] = 83
              "01010100" when "11001111", -- t[207] = 84
              "01010101" when "11010000", -- t[208] = 85
              "01010101" when "11010001", -- t[209] = 85
              "01010110" when "11010010", -- t[210] = 86
              "01010111" when "11010011", -- t[211] = 87
              "01011000" when "11010100", -- t[212] = 88
              "01011001" when "11010101", -- t[213] = 89
              "01011010" when "11010110", -- t[214] = 90
              "01011010" when "11010111", -- t[215] = 90
              "01011011" when "11011000", -- t[216] = 91
              "01011100" when "11011001", -- t[217] = 92
              "01011101" when "11011010", -- t[218] = 93
              "01011110" when "11011011", -- t[219] = 94
              "01011111" when "11011100", -- t[220] = 95
              "01100000" when "11011101", -- t[221] = 96
              "01100000" when "11011110", -- t[222] = 96
              "01100001" when "11011111", -- t[223] = 97
              "01100010" when "11100000", -- t[224] = 98
              "01100011" when "11100001", -- t[225] = 99
              "01100100" when "11100010", -- t[226] = 100
              "01100101" when "11100011", -- t[227] = 101
              "01100110" when "11100100", -- t[228] = 102
              "01100111" when "11100101", -- t[229] = 103
              "01101000" when "11100110", -- t[230] = 104
              "01101000" when "11100111", -- t[231] = 104
              "01101001" when "11101000", -- t[232] = 105
              "01101010" when "11101001", -- t[233] = 106
              "01101011" when "11101010", -- t[234] = 107
              "01101100" when "11101011", -- t[235] = 108
              "01101101" when "11101100", -- t[236] = 109
              "01101110" when "11101101", -- t[237] = 110
              "01101111" when "11101110", -- t[238] = 111
              "01110000" when "11101111", -- t[239] = 112
              "01110001" when "11110000", -- t[240] = 113
              "01110010" when "11110001", -- t[241] = 114
              "01110011" when "11110010", -- t[242] = 115
              "01110100" when "11110011", -- t[243] = 116
              "01110101" when "11110100", -- t[244] = 117
              "01110110" when "11110101", -- t[245] = 118
              "01110110" when "11110110", -- t[246] = 118
              "01110111" when "11110111", -- t[247] = 119
              "01111000" when "11111000", -- t[248] = 120
              "01111001" when "11111001", -- t[249] = 121
              "01111010" when "11111010", -- t[250] = 122
              "01111011" when "11111011", -- t[251] = 123
              "01111100" when "11111100", -- t[252] = 124
              "01111101" when "11111101", -- t[253] = 125
              "01111110" when "11111110", -- t[254] = 126
              "01111111" when "11111111", -- t[255] = 127
              "--------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_18 is
  port ( nY2    : in  std_logic_vector(6 downto 0);
         nExpY2 : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_18 is
begin

  with nY2 select
    nExpY2 <= "0000000" when "0000000", -- t[0] = 0
              "0000000" when "0000001", -- t[1] = 0
              "0000000" when "0000010", -- t[2] = 0
              "0000000" when "0000011", -- t[3] = 0
              "0000000" when "0000100", -- t[4] = 0
              "0000000" when "0000101", -- t[5] = 0
              "0000000" when "0000110", -- t[6] = 0
              "0000000" when "0000111", -- t[7] = 0
              "0000000" when "0001000", -- t[8] = 0
              "0000000" when "0001001", -- t[9] = 0
              "0000000" when "0001010", -- t[10] = 0
              "0000000" when "0001011", -- t[11] = 0
              "0000001" when "0001100", -- t[12] = 1
              "0000001" when "0001101", -- t[13] = 1
              "0000001" when "0001110", -- t[14] = 1
              "0000001" when "0001111", -- t[15] = 1
              "0000001" when "0010000", -- t[16] = 1
              "0000001" when "0010001", -- t[17] = 1
              "0000001" when "0010010", -- t[18] = 1
              "0000001" when "0010011", -- t[19] = 1
              "0000010" when "0010100", -- t[20] = 2
              "0000010" when "0010101", -- t[21] = 2
              "0000010" when "0010110", -- t[22] = 2
              "0000010" when "0010111", -- t[23] = 2
              "0000010" when "0011000", -- t[24] = 2
              "0000010" when "0011001", -- t[25] = 2
              "0000011" when "0011010", -- t[26] = 3
              "0000011" when "0011011", -- t[27] = 3
              "0000011" when "0011100", -- t[28] = 3
              "0000011" when "0011101", -- t[29] = 3
              "0000100" when "0011110", -- t[30] = 4
              "0000100" when "0011111", -- t[31] = 4
              "0000100" when "0100000", -- t[32] = 4
              "0000100" when "0100001", -- t[33] = 4
              "0000101" when "0100010", -- t[34] = 5
              "0000101" when "0100011", -- t[35] = 5
              "0000101" when "0100100", -- t[36] = 5
              "0000101" when "0100101", -- t[37] = 5
              "0000110" when "0100110", -- t[38] = 6
              "0000110" when "0100111", -- t[39] = 6
              "0000110" when "0101000", -- t[40] = 6
              "0000111" when "0101001", -- t[41] = 7
              "0000111" when "0101010", -- t[42] = 7
              "0000111" when "0101011", -- t[43] = 7
              "0001000" when "0101100", -- t[44] = 8
              "0001000" when "0101101", -- t[45] = 8
              "0001000" when "0101110", -- t[46] = 8
              "0001001" when "0101111", -- t[47] = 9
              "0001001" when "0110000", -- t[48] = 9
              "0001001" when "0110001", -- t[49] = 9
              "0001010" when "0110010", -- t[50] = 10
              "0001010" when "0110011", -- t[51] = 10
              "0001011" when "0110100", -- t[52] = 11
              "0001011" when "0110101", -- t[53] = 11
              "0001011" when "0110110", -- t[54] = 11
              "0001100" when "0110111", -- t[55] = 12
              "0001100" when "0111000", -- t[56] = 12
              "0001101" when "0111001", -- t[57] = 13
              "0001101" when "0111010", -- t[58] = 13
              "0001110" when "0111011", -- t[59] = 14
              "0001110" when "0111100", -- t[60] = 14
              "0001111" when "0111101", -- t[61] = 15
              "0001111" when "0111110", -- t[62] = 15
              "0010000" when "0111111", -- t[63] = 16
              "0010000" when "1000000", -- t[64] = 16
              "0010001" when "1000001", -- t[65] = 17
              "0010001" when "1000010", -- t[66] = 17
              "0010010" when "1000011", -- t[67] = 18
              "0010010" when "1000100", -- t[68] = 18
              "0010011" when "1000101", -- t[69] = 19
              "0010011" when "1000110", -- t[70] = 19
              "0010100" when "1000111", -- t[71] = 20
              "0010100" when "1001000", -- t[72] = 20
              "0010101" when "1001001", -- t[73] = 21
              "0010101" when "1001010", -- t[74] = 21
              "0010110" when "1001011", -- t[75] = 22
              "0010111" when "1001100", -- t[76] = 23
              "0010111" when "1001101", -- t[77] = 23
              "0011000" when "1001110", -- t[78] = 24
              "0011000" when "1001111", -- t[79] = 24
              "0011001" when "1010000", -- t[80] = 25
              "0011010" when "1010001", -- t[81] = 26
              "0011010" when "1010010", -- t[82] = 26
              "0011011" when "1010011", -- t[83] = 27
              "0011100" when "1010100", -- t[84] = 28
              "0011100" when "1010101", -- t[85] = 28
              "0011101" when "1010110", -- t[86] = 29
              "0011110" when "1010111", -- t[87] = 30
              "0011110" when "1011000", -- t[88] = 30
              "0011111" when "1011001", -- t[89] = 31
              "0100000" when "1011010", -- t[90] = 32
              "0100000" when "1011011", -- t[91] = 32
              "0100001" when "1011100", -- t[92] = 33
              "0100010" when "1011101", -- t[93] = 34
              "0100011" when "1011110", -- t[94] = 35
              "0100011" when "1011111", -- t[95] = 35
              "0100100" when "1100000", -- t[96] = 36
              "0100101" when "1100001", -- t[97] = 37
              "0100110" when "1100010", -- t[98] = 38
              "0100110" when "1100011", -- t[99] = 38
              "0100111" when "1100100", -- t[100] = 39
              "0101000" when "1100101", -- t[101] = 40
              "0101001" when "1100110", -- t[102] = 41
              "0101001" when "1100111", -- t[103] = 41
              "0101010" when "1101000", -- t[104] = 42
              "0101011" when "1101001", -- t[105] = 43
              "0101100" when "1101010", -- t[106] = 44
              "0101101" when "1101011", -- t[107] = 45
              "0101110" when "1101100", -- t[108] = 46
              "0101110" when "1101101", -- t[109] = 46
              "0101111" when "1101110", -- t[110] = 47
              "0110000" when "1101111", -- t[111] = 48
              "0110001" when "1110000", -- t[112] = 49
              "0110010" when "1110001", -- t[113] = 50
              "0110011" when "1110010", -- t[114] = 51
              "0110100" when "1110011", -- t[115] = 52
              "0110101" when "1110100", -- t[116] = 53
              "0110110" when "1110101", -- t[117] = 54
              "0110110" when "1110110", -- t[118] = 54
              "0110111" when "1110111", -- t[119] = 55
              "0111000" when "1111000", -- t[120] = 56
              "0111001" when "1111001", -- t[121] = 57
              "0111010" when "1111010", -- t[122] = 58
              "0111011" when "1111011", -- t[123] = 59
              "0111100" when "1111100", -- t[124] = 60
              "0111101" when "1111101", -- t[125] = 61
              "0111110" when "1111110", -- t[126] = 62
              "0111111" when "1111111", -- t[127] = 63
              "-------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_19 is
  port ( nY2    : in  std_logic_vector(7 downto 0);
         nExpY2 : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_19 is
begin

  with nY2 select
    nExpY2 <= "00000000" when "00000000", -- t[0] = 0
              "00000000" when "00000001", -- t[1] = 0
              "00000000" when "00000010", -- t[2] = 0
              "00000000" when "00000011", -- t[3] = 0
              "00000000" when "00000100", -- t[4] = 0
              "00000000" when "00000101", -- t[5] = 0
              "00000000" when "00000110", -- t[6] = 0
              "00000000" when "00000111", -- t[7] = 0
              "00000000" when "00001000", -- t[8] = 0
              "00000000" when "00001001", -- t[9] = 0
              "00000000" when "00001010", -- t[10] = 0
              "00000000" when "00001011", -- t[11] = 0
              "00000000" when "00001100", -- t[12] = 0
              "00000000" when "00001101", -- t[13] = 0
              "00000000" when "00001110", -- t[14] = 0
              "00000000" when "00001111", -- t[15] = 0
              "00000001" when "00010000", -- t[16] = 1
              "00000001" when "00010001", -- t[17] = 1
              "00000001" when "00010010", -- t[18] = 1
              "00000001" when "00010011", -- t[19] = 1
              "00000001" when "00010100", -- t[20] = 1
              "00000001" when "00010101", -- t[21] = 1
              "00000001" when "00010110", -- t[22] = 1
              "00000001" when "00010111", -- t[23] = 1
              "00000001" when "00011000", -- t[24] = 1
              "00000001" when "00011001", -- t[25] = 1
              "00000001" when "00011010", -- t[26] = 1
              "00000001" when "00011011", -- t[27] = 1
              "00000010" when "00011100", -- t[28] = 2
              "00000010" when "00011101", -- t[29] = 2
              "00000010" when "00011110", -- t[30] = 2
              "00000010" when "00011111", -- t[31] = 2
              "00000010" when "00100000", -- t[32] = 2
              "00000010" when "00100001", -- t[33] = 2
              "00000010" when "00100010", -- t[34] = 2
              "00000010" when "00100011", -- t[35] = 2
              "00000011" when "00100100", -- t[36] = 3
              "00000011" when "00100101", -- t[37] = 3
              "00000011" when "00100110", -- t[38] = 3
              "00000011" when "00100111", -- t[39] = 3
              "00000011" when "00101000", -- t[40] = 3
              "00000011" when "00101001", -- t[41] = 3
              "00000011" when "00101010", -- t[42] = 3
              "00000100" when "00101011", -- t[43] = 4
              "00000100" when "00101100", -- t[44] = 4
              "00000100" when "00101101", -- t[45] = 4
              "00000100" when "00101110", -- t[46] = 4
              "00000100" when "00101111", -- t[47] = 4
              "00000101" when "00110000", -- t[48] = 5
              "00000101" when "00110001", -- t[49] = 5
              "00000101" when "00110010", -- t[50] = 5
              "00000101" when "00110011", -- t[51] = 5
              "00000101" when "00110100", -- t[52] = 5
              "00000101" when "00110101", -- t[53] = 5
              "00000110" when "00110110", -- t[54] = 6
              "00000110" when "00110111", -- t[55] = 6
              "00000110" when "00111000", -- t[56] = 6
              "00000110" when "00111001", -- t[57] = 6
              "00000111" when "00111010", -- t[58] = 7
              "00000111" when "00111011", -- t[59] = 7
              "00000111" when "00111100", -- t[60] = 7
              "00000111" when "00111101", -- t[61] = 7
              "00001000" when "00111110", -- t[62] = 8
              "00001000" when "00111111", -- t[63] = 8
              "00001000" when "01000000", -- t[64] = 8
              "00001000" when "01000001", -- t[65] = 8
              "00001001" when "01000010", -- t[66] = 9
              "00001001" when "01000011", -- t[67] = 9
              "00001001" when "01000100", -- t[68] = 9
              "00001001" when "01000101", -- t[69] = 9
              "00001010" when "01000110", -- t[70] = 10
              "00001010" when "01000111", -- t[71] = 10
              "00001010" when "01001000", -- t[72] = 10
              "00001010" when "01001001", -- t[73] = 10
              "00001011" when "01001010", -- t[74] = 11
              "00001011" when "01001011", -- t[75] = 11
              "00001011" when "01001100", -- t[76] = 11
              "00001100" when "01001101", -- t[77] = 12
              "00001100" when "01001110", -- t[78] = 12
              "00001100" when "01001111", -- t[79] = 12
              "00001101" when "01010000", -- t[80] = 13
              "00001101" when "01010001", -- t[81] = 13
              "00001101" when "01010010", -- t[82] = 13
              "00001101" when "01010011", -- t[83] = 13
              "00001110" when "01010100", -- t[84] = 14
              "00001110" when "01010101", -- t[85] = 14
              "00001110" when "01010110", -- t[86] = 14
              "00001111" when "01010111", -- t[87] = 15
              "00001111" when "01011000", -- t[88] = 15
              "00001111" when "01011001", -- t[89] = 15
              "00010000" when "01011010", -- t[90] = 16
              "00010000" when "01011011", -- t[91] = 16
              "00010001" when "01011100", -- t[92] = 17
              "00010001" when "01011101", -- t[93] = 17
              "00010001" when "01011110", -- t[94] = 17
              "00010010" when "01011111", -- t[95] = 18
              "00010010" when "01100000", -- t[96] = 18
              "00010010" when "01100001", -- t[97] = 18
              "00010011" when "01100010", -- t[98] = 19
              "00010011" when "01100011", -- t[99] = 19
              "00010100" when "01100100", -- t[100] = 20
              "00010100" when "01100101", -- t[101] = 20
              "00010100" when "01100110", -- t[102] = 20
              "00010101" when "01100111", -- t[103] = 21
              "00010101" when "01101000", -- t[104] = 21
              "00010110" when "01101001", -- t[105] = 22
              "00010110" when "01101010", -- t[106] = 22
              "00010110" when "01101011", -- t[107] = 22
              "00010111" when "01101100", -- t[108] = 23
              "00010111" when "01101101", -- t[109] = 23
              "00011000" when "01101110", -- t[110] = 24
              "00011000" when "01101111", -- t[111] = 24
              "00011001" when "01110000", -- t[112] = 25
              "00011001" when "01110001", -- t[113] = 25
              "00011001" when "01110010", -- t[114] = 25
              "00011010" when "01110011", -- t[115] = 26
              "00011010" when "01110100", -- t[116] = 26
              "00011011" when "01110101", -- t[117] = 27
              "00011011" when "01110110", -- t[118] = 27
              "00011100" when "01110111", -- t[119] = 28
              "00011100" when "01111000", -- t[120] = 28
              "00011101" when "01111001", -- t[121] = 29
              "00011101" when "01111010", -- t[122] = 29
              "00011110" when "01111011", -- t[123] = 30
              "00011110" when "01111100", -- t[124] = 30
              "00011111" when "01111101", -- t[125] = 31
              "00011111" when "01111110", -- t[126] = 31
              "00100000" when "01111111", -- t[127] = 32
              "00100000" when "10000000", -- t[128] = 32
              "00100001" when "10000001", -- t[129] = 33
              "00100001" when "10000010", -- t[130] = 33
              "00100010" when "10000011", -- t[131] = 34
              "00100010" when "10000100", -- t[132] = 34
              "00100011" when "10000101", -- t[133] = 35
              "00100011" when "10000110", -- t[134] = 35
              "00100100" when "10000111", -- t[135] = 36
              "00100100" when "10001000", -- t[136] = 36
              "00100101" when "10001001", -- t[137] = 37
              "00100101" when "10001010", -- t[138] = 37
              "00100110" when "10001011", -- t[139] = 38
              "00100110" when "10001100", -- t[140] = 38
              "00100111" when "10001101", -- t[141] = 39
              "00100111" when "10001110", -- t[142] = 39
              "00101000" when "10001111", -- t[143] = 40
              "00101001" when "10010000", -- t[144] = 41
              "00101001" when "10010001", -- t[145] = 41
              "00101010" when "10010010", -- t[146] = 42
              "00101010" when "10010011", -- t[147] = 42
              "00101011" when "10010100", -- t[148] = 43
              "00101011" when "10010101", -- t[149] = 43
              "00101100" when "10010110", -- t[150] = 44
              "00101101" when "10010111", -- t[151] = 45
              "00101101" when "10011000", -- t[152] = 45
              "00101110" when "10011001", -- t[153] = 46
              "00101110" when "10011010", -- t[154] = 46
              "00101111" when "10011011", -- t[155] = 47
              "00110000" when "10011100", -- t[156] = 48
              "00110000" when "10011101", -- t[157] = 48
              "00110001" when "10011110", -- t[158] = 49
              "00110001" when "10011111", -- t[159] = 49
              "00110010" when "10100000", -- t[160] = 50
              "00110011" when "10100001", -- t[161] = 51
              "00110011" when "10100010", -- t[162] = 51
              "00110100" when "10100011", -- t[163] = 52
              "00110101" when "10100100", -- t[164] = 53
              "00110101" when "10100101", -- t[165] = 53
              "00110110" when "10100110", -- t[166] = 54
              "00110111" when "10100111", -- t[167] = 55
              "00110111" when "10101000", -- t[168] = 55
              "00111000" when "10101001", -- t[169] = 56
              "00111000" when "10101010", -- t[170] = 56
              "00111001" when "10101011", -- t[171] = 57
              "00111010" when "10101100", -- t[172] = 58
              "00111011" when "10101101", -- t[173] = 59
              "00111011" when "10101110", -- t[174] = 59
              "00111100" when "10101111", -- t[175] = 60
              "00111101" when "10110000", -- t[176] = 61
              "00111101" when "10110001", -- t[177] = 61
              "00111110" when "10110010", -- t[178] = 62
              "00111111" when "10110011", -- t[179] = 63
              "00111111" when "10110100", -- t[180] = 63
              "01000000" when "10110101", -- t[181] = 64
              "01000001" when "10110110", -- t[182] = 65
              "01000001" when "10110111", -- t[183] = 65
              "01000010" when "10111000", -- t[184] = 66
              "01000011" when "10111001", -- t[185] = 67
              "01000100" when "10111010", -- t[186] = 68
              "01000100" when "10111011", -- t[187] = 68
              "01000101" when "10111100", -- t[188] = 69
              "01000110" when "10111101", -- t[189] = 70
              "01000111" when "10111110", -- t[190] = 71
              "01000111" when "10111111", -- t[191] = 71
              "01001000" when "11000000", -- t[192] = 72
              "01001001" when "11000001", -- t[193] = 73
              "01001010" when "11000010", -- t[194] = 74
              "01001010" when "11000011", -- t[195] = 74
              "01001011" when "11000100", -- t[196] = 75
              "01001100" when "11000101", -- t[197] = 76
              "01001101" when "11000110", -- t[198] = 77
              "01001101" when "11000111", -- t[199] = 77
              "01001110" when "11001000", -- t[200] = 78
              "01001111" when "11001001", -- t[201] = 79
              "01010000" when "11001010", -- t[202] = 80
              "01010001" when "11001011", -- t[203] = 81
              "01010001" when "11001100", -- t[204] = 81
              "01010010" when "11001101", -- t[205] = 82
              "01010011" when "11001110", -- t[206] = 83
              "01010100" when "11001111", -- t[207] = 84
              "01010101" when "11010000", -- t[208] = 85
              "01010101" when "11010001", -- t[209] = 85
              "01010110" when "11010010", -- t[210] = 86
              "01010111" when "11010011", -- t[211] = 87
              "01011000" when "11010100", -- t[212] = 88
              "01011001" when "11010101", -- t[213] = 89
              "01011010" when "11010110", -- t[214] = 90
              "01011010" when "11010111", -- t[215] = 90
              "01011011" when "11011000", -- t[216] = 91
              "01011100" when "11011001", -- t[217] = 92
              "01011101" when "11011010", -- t[218] = 93
              "01011110" when "11011011", -- t[219] = 94
              "01011111" when "11011100", -- t[220] = 95
              "01011111" when "11011101", -- t[221] = 95
              "01100000" when "11011110", -- t[222] = 96
              "01100001" when "11011111", -- t[223] = 97
              "01100010" when "11100000", -- t[224] = 98
              "01100011" when "11100001", -- t[225] = 99
              "01100100" when "11100010", -- t[226] = 100
              "01100101" when "11100011", -- t[227] = 101
              "01100110" when "11100100", -- t[228] = 102
              "01100111" when "11100101", -- t[229] = 103
              "01100111" when "11100110", -- t[230] = 103
              "01101000" when "11100111", -- t[231] = 104
              "01101001" when "11101000", -- t[232] = 105
              "01101010" when "11101001", -- t[233] = 106
              "01101011" when "11101010", -- t[234] = 107
              "01101100" when "11101011", -- t[235] = 108
              "01101101" when "11101100", -- t[236] = 109
              "01101110" when "11101101", -- t[237] = 110
              "01101111" when "11101110", -- t[238] = 111
              "01110000" when "11101111", -- t[239] = 112
              "01110001" when "11110000", -- t[240] = 113
              "01110010" when "11110001", -- t[241] = 114
              "01110011" when "11110010", -- t[242] = 115
              "01110011" when "11110011", -- t[243] = 115
              "01110100" when "11110100", -- t[244] = 116
              "01110101" when "11110101", -- t[245] = 117
              "01110110" when "11110110", -- t[246] = 118
              "01110111" when "11110111", -- t[247] = 119
              "01111000" when "11111000", -- t[248] = 120
              "01111001" when "11111001", -- t[249] = 121
              "01111010" when "11111010", -- t[250] = 122
              "01111011" when "11111011", -- t[251] = 123
              "01111100" when "11111100", -- t[252] = 124
              "01111101" when "11111101", -- t[253] = 125
              "01111110" when "11111110", -- t[254] = 126
              "01111111" when "11111111", -- t[255] = 127
              "--------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function e^x-x-1.
-- wI = 9; wO = 9.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 5; beta = 4;
--   T_0 (ROM):     alpha_0 = 5; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 4; beta_1 = 4.
-- Guard bits: g = 1.
-- Command line: exp 9 9 1   rom 5 0   pm 4 4  ah 4 4 4  0 1  4 4 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 5; beta_0 = 0; wO_0 = 10.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_20_t0 is
  port ( a : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_20_t0 is
  signal x0   : std_logic_vector(4 downto 0);
  signal r0   : std_logic_vector(9 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "0000000001" when "00000", -- t[0] = 1
          "0000000011" when "00001", -- t[1] = 3
          "0000000111" when "00010", -- t[2] = 7
          "0000001101" when "00011", -- t[3] = 13
          "0000010101" when "00100", -- t[4] = 21
          "0000011111" when "00101", -- t[5] = 31
          "0000101011" when "00110", -- t[6] = 43
          "0000111001" when "00111", -- t[7] = 57
          "0001001001" when "01000", -- t[8] = 73
          "0001011011" when "01001", -- t[9] = 91
          "0001101111" when "01010", -- t[10] = 111
          "0010000101" when "01011", -- t[11] = 133
          "0010011101" when "01100", -- t[12] = 157
          "0010110111" when "01101", -- t[13] = 183
          "0011010011" when "01110", -- t[14] = 211
          "0011110000" when "01111", -- t[15] = 240
          "0100010000" when "10000", -- t[16] = 272
          "0100110010" when "10001", -- t[17] = 306
          "0101010110" when "10010", -- t[18] = 342
          "0101111100" when "10011", -- t[19] = 380
          "0110100100" when "10100", -- t[20] = 420
          "0111001110" when "10101", -- t[21] = 462
          "0111111010" when "10110", -- t[22] = 506
          "1000101000" when "10111", -- t[23] = 552
          "1001011000" when "11000", -- t[24] = 600
          "1010001010" when "11001", -- t[25] = 650
          "1010111110" when "11010", -- t[26] = 702
          "1011110100" when "11011", -- t[27] = 756
          "1100101100" when "11100", -- t[28] = 812
          "1101100110" when "11101", -- t[29] = 870
          "1110100010" when "11110", -- t[30] = 930
          "1111100000" when "11111", -- t[31] = 992
          "----------" when others;

  r(9 downto 0) <= r0;
  r(10 downto 10) <= (10 downto 10 => ('0'));
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 4; mu_1 = 4; lambda_1 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_20_t1_pow is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_20_t1_pow is
  signal pp0 : std_logic_vector(2 downto 0);
  signal r0 : std_logic_vector(2 downto 0);
begin
  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(2 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 4; sigma'_1,1 = 3; wO_1,1 = 5.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_20_t1_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         s : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_20_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a & s;

  with x select
    r <= "00000" when "0000000", -- t[0] = 0
         "00000" when "0000001", -- t[1] = 0
         "00000" when "0000010", -- t[2] = 0
         "00000" when "0000011", -- t[3] = 0
         "00000" when "0000100", -- t[4] = 0
         "00000" when "0000101", -- t[5] = 0
         "00000" when "0000110", -- t[6] = 0
         "00000" when "0000111", -- t[7] = 0
         "00000" when "0001000", -- t[8] = 0
         "00000" when "0001001", -- t[9] = 0
         "00000" when "0001010", -- t[10] = 0
         "00001" when "0001011", -- t[11] = 1
         "00001" when "0001100", -- t[12] = 1
         "00010" when "0001101", -- t[13] = 2
         "00010" when "0001110", -- t[14] = 2
         "00010" when "0001111", -- t[15] = 2
         "00000" when "0010000", -- t[16] = 0
         "00000" when "0010001", -- t[17] = 0
         "00001" when "0010010", -- t[18] = 1
         "00010" when "0010011", -- t[19] = 2
         "00010" when "0010100", -- t[20] = 2
         "00011" when "0010101", -- t[21] = 3
         "00100" when "0010110", -- t[22] = 4
         "00100" when "0010111", -- t[23] = 4
         "00000" when "0011000", -- t[24] = 0
         "00001" when "0011001", -- t[25] = 1
         "00010" when "0011010", -- t[26] = 2
         "00011" when "0011011", -- t[27] = 3
         "00011" when "0011100", -- t[28] = 3
         "00100" when "0011101", -- t[29] = 4
         "00101" when "0011110", -- t[30] = 5
         "00110" when "0011111", -- t[31] = 6
         "00000" when "0100000", -- t[32] = 0
         "00001" when "0100001", -- t[33] = 1
         "00010" when "0100010", -- t[34] = 2
         "00011" when "0100011", -- t[35] = 3
         "00101" when "0100100", -- t[36] = 5
         "00110" when "0100101", -- t[37] = 6
         "00111" when "0100110", -- t[38] = 7
         "01000" when "0100111", -- t[39] = 8
         "00000" when "0101000", -- t[40] = 0
         "00010" when "0101001", -- t[41] = 2
         "00011" when "0101010", -- t[42] = 3
         "00100" when "0101011", -- t[43] = 4
         "00110" when "0101100", -- t[44] = 6
         "00111" when "0101101", -- t[45] = 7
         "01000" when "0101110", -- t[46] = 8
         "01010" when "0101111", -- t[47] = 10
         "00000" when "0110000", -- t[48] = 0
         "00010" when "0110001", -- t[49] = 2
         "00100" when "0110010", -- t[50] = 4
         "00101" when "0110011", -- t[51] = 5
         "00111" when "0110100", -- t[52] = 7
         "01000" when "0110101", -- t[53] = 8
         "01010" when "0110110", -- t[54] = 10
         "01100" when "0110111", -- t[55] = 12
         "00000" when "0111000", -- t[56] = 0
         "00010" when "0111001", -- t[57] = 2
         "00100" when "0111010", -- t[58] = 4
         "00110" when "0111011", -- t[59] = 6
         "01000" when "0111100", -- t[60] = 8
         "01010" when "0111101", -- t[61] = 10
         "01100" when "0111110", -- t[62] = 12
         "01110" when "0111111", -- t[63] = 14
         "00001" when "1000000", -- t[64] = 1
         "00011" when "1000001", -- t[65] = 3
         "00101" when "1000010", -- t[66] = 5
         "00111" when "1000011", -- t[67] = 7
         "01001" when "1000100", -- t[68] = 9
         "01011" when "1000101", -- t[69] = 11
         "01101" when "1000110", -- t[70] = 13
         "01111" when "1000111", -- t[71] = 15
         "00001" when "1001000", -- t[72] = 1
         "00011" when "1001001", -- t[73] = 3
         "00101" when "1001010", -- t[74] = 5
         "01000" when "1001011", -- t[75] = 8
         "01010" when "1001100", -- t[76] = 10
         "01101" when "1001101", -- t[77] = 13
         "01111" when "1001110", -- t[78] = 15
         "10001" when "1001111", -- t[79] = 17
         "00001" when "1010000", -- t[80] = 1
         "00011" when "1010001", -- t[81] = 3
         "00110" when "1010010", -- t[82] = 6
         "01001" when "1010011", -- t[83] = 9
         "01011" when "1010100", -- t[84] = 11
         "01110" when "1010101", -- t[85] = 14
         "10001" when "1010110", -- t[86] = 17
         "10011" when "1010111", -- t[87] = 19
         "00001" when "1011000", -- t[88] = 1
         "00100" when "1011001", -- t[89] = 4
         "00111" when "1011010", -- t[90] = 7
         "01010" when "1011011", -- t[91] = 10
         "01100" when "1011100", -- t[92] = 12
         "01111" when "1011101", -- t[93] = 15
         "10010" when "1011110", -- t[94] = 18
         "10101" when "1011111", -- t[95] = 21
         "00001" when "1100000", -- t[96] = 1
         "00100" when "1100001", -- t[97] = 4
         "00111" when "1100010", -- t[98] = 7
         "01010" when "1100011", -- t[99] = 10
         "01110" when "1100100", -- t[100] = 14
         "10001" when "1100101", -- t[101] = 17
         "10100" when "1100110", -- t[102] = 20
         "10111" when "1100111", -- t[103] = 23
         "00001" when "1101000", -- t[104] = 1
         "00101" when "1101001", -- t[105] = 5
         "01000" when "1101010", -- t[106] = 8
         "01011" when "1101011", -- t[107] = 11
         "01111" when "1101100", -- t[108] = 15
         "10010" when "1101101", -- t[109] = 18
         "10101" when "1101110", -- t[110] = 21
         "11001" when "1101111", -- t[111] = 25
         "00001" when "1110000", -- t[112] = 1
         "00101" when "1110001", -- t[113] = 5
         "01001" when "1110010", -- t[114] = 9
         "01100" when "1110011", -- t[115] = 12
         "10000" when "1110100", -- t[116] = 16
         "10011" when "1110101", -- t[117] = 19
         "10111" when "1110110", -- t[118] = 23
         "11011" when "1110111", -- t[119] = 27
         "00001" when "1111000", -- t[120] = 1
         "00101" when "1111001", -- t[121] = 5
         "01001" when "1111010", -- t[122] = 9
         "01101" when "1111011", -- t[123] = 13
         "10001" when "1111100", -- t[124] = 17
         "10101" when "1111101", -- t[125] = 21
         "11001" when "1111110", -- t[126] = 25
         "11101" when "1111111", -- t[127] = 29
         "-----" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 4; beta_1 = 4; lambda_1 = 4;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (ROM):  alpha_1,1 = 4; rho_1,1 = 0; sigma_1,1 = 4; wO_1,1 = 5.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_20_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_20_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(2 downto 0);
  signal s      : std_logic_vector(3 downto 0);
  component fp_exp_exp_y2_20_t1_pow is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  signal a_1    : std_logic_vector(3 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(2 downto 0);
  signal r0_1   : std_logic_vector(4 downto 0);
  signal r_1    : std_logic_vector(10 downto 0);
  component fp_exp_exp_y2_20_t1_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;
begin
  sign <= not b(3);
  b0 <= b(2 downto 0) xor (2 downto 0 => sign);

  pow : fp_exp_exp_y2_20_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(3 downto 0);
  sign_1 <= not s(3);
  s_1 <= s(2 downto 0) xor (2 downto 0 => sign_1);
  t_1 : fp_exp_exp_y2_20_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_1 );
  r_1(4 downto 0) <=
    r0_1 xor (4 downto 0 => ((sign xor sign_1)));
  r_1(10 downto 5) <= (10 downto 5 => ((sign xor sign_1)));

  r <= r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_20_t1_clk is
  port ( a   : in  std_logic_vector(3 downto 0);
         b   : in  std_logic_vector(3 downto 0);
         r   : out std_logic_vector(10 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_20_t1_clk is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(2 downto 0);
  signal s      : std_logic_vector(3 downto 0);
  component fp_exp_exp_y2_20_t1_pow is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  signal a_1     : std_logic_vector(3 downto 0);
  signal sign_1  : std_logic;
  signal s_1     : std_logic_vector(2 downto 0);
  signal r0_10   : std_logic_vector(4 downto 0);
  signal r0_1r   : std_logic_vector(4 downto 0);
  signal r_1     : std_logic_vector(10 downto 0);
  signal sign_10 : std_logic;
  signal sign_1r : std_logic;
  component fp_exp_exp_y2_20_t1_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;
begin
  sign <= not b(3);
  b0 <= b(2 downto 0) xor (2 downto 0 => sign);

  pow : fp_exp_exp_y2_20_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(3 downto 0);
  sign_1 <= not s(3);
  s_1 <= s(2 downto 0) xor (2 downto 0 => sign_1);
  sign_10 <= sign xor sign_1;
  t_1 : fp_exp_exp_y2_20_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_10 );
  r_1(4 downto 0) <=
    r0_1r xor (4 downto 0 => sign_1r);
  r_1(10 downto 5) <= (10 downto 5 => sign_1r);

  process(clk)
  begin
    if clk'event and clk = '1' then
      r0_1r   <= r0_10;
      sign_1r <= sign_10;
    end if;
  end process;

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_20 is
  port ( x : in  std_logic_vector(8 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_20 is
  signal a_0 : std_logic_vector(4 downto 0);
  signal r_0 : std_logic_vector(10 downto 0);
  component fp_exp_exp_y2_20_t0 is
    port ( a : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  signal a_1 : std_logic_vector(3 downto 0);
  signal b_1 : std_logic_vector(3 downto 0);
  signal r_1 : std_logic_vector(10 downto 0);
  component fp_exp_exp_y2_20_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  signal sum : std_logic_vector(10 downto 0);
begin
  a_0 <= x(8 downto 4);
  t_0 : fp_exp_exp_y2_20_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(8 downto 5);
  b_1 <= x(3 downto 0);
  t_1 : fp_exp_exp_y2_20_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  sum <= r_0 + r_1;
  r <= sum(10 downto 1);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_20_clk is
  port ( x   : in  std_logic_vector(8 downto 0);
         r   : out std_logic_vector(9 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_20_clk is
  signal a_x0 : std_logic_vector(4 downto 0);
  signal a_xr : std_logic_vector(4 downto 0);
  signal r_0  : std_logic_vector(10 downto 0);
  component fp_exp_exp_y2_20_t0 is
    port ( a : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  signal a_1 : std_logic_vector(3 downto 0);
  signal b_1 : std_logic_vector(3 downto 0);
  signal r_1 : std_logic_vector(10 downto 0);
  component fp_exp_exp_y2_20_t1_clk is
    port ( a   : in  std_logic_vector(3 downto 0);
           b   : in  std_logic_vector(3 downto 0);
           r   : out std_logic_vector(10 downto 0);
           clk : in  std_logic );
  end component;

  signal sum : std_logic_vector(10 downto 0);
begin
  a_x0 <= x(8 downto 4);
  t_0 : fp_exp_exp_y2_20_t0
    port map ( a => a_xr,
               r => r_0 );

  process(clk)
  begin
    if clk'event and clk = '1' then
      a_xr <= a_x0;
    end if;
  end process;

  a_1 <= x(8 downto 5);
  b_1 <= x(3 downto 0);
  t_1 : fp_exp_exp_y2_20_t1_clk
    port map ( a   => a_1,
               b   => b_1,
               r   => r_1,
               clk => clk );

  sum <= r_0 + r_1;
  r <= sum(10 downto 1);
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function e^x-x-1.
-- wI = 10; wO = 10.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 6; beta = 4;
--   T_0 (ROM):     alpha_0 = 6; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 4; beta_1 = 4.
-- Guard bits: g = 2.
-- Command line: exp 10 10 1   rom 6 0   pm 4 4  ah 4 4 4  0 1  4 4 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 6; beta_0 = 0; wO_0 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_21_t0 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_21_t0 is
  signal x0   : std_logic_vector(5 downto 0);
  signal r0   : std_logic_vector(11 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "000000000010" when "000000", -- t[0] = 2
          "000000000100" when "000001", -- t[1] = 4
          "000000001000" when "000010", -- t[2] = 8
          "000000001110" when "000011", -- t[3] = 14
          "000000010110" when "000100", -- t[4] = 22
          "000000100000" when "000101", -- t[5] = 32
          "000000101100" when "000110", -- t[6] = 44
          "000000111010" when "000111", -- t[7] = 58
          "000001001010" when "001000", -- t[8] = 74
          "000001011100" when "001001", -- t[9] = 92
          "000001110000" when "001010", -- t[10] = 112
          "000010000110" when "001011", -- t[11] = 134
          "000010011110" when "001100", -- t[12] = 158
          "000010111000" when "001101", -- t[13] = 184
          "000011010011" when "001110", -- t[14] = 211
          "000011110001" when "001111", -- t[15] = 241
          "000100010001" when "010000", -- t[16] = 273
          "000100110011" when "010001", -- t[17] = 307
          "000101010111" when "010010", -- t[18] = 343
          "000101111101" when "010011", -- t[19] = 381
          "000110100101" when "010100", -- t[20] = 421
          "000111001111" when "010101", -- t[21] = 463
          "000111111011" when "010110", -- t[22] = 507
          "001000101001" when "010111", -- t[23] = 553
          "001001011001" when "011000", -- t[24] = 601
          "001010001011" when "011001", -- t[25] = 651
          "001010111111" when "011010", -- t[26] = 703
          "001011110101" when "011011", -- t[27] = 757
          "001100101101" when "011100", -- t[28] = 813
          "001101100111" when "011101", -- t[29] = 871
          "001110100011" when "011110", -- t[30] = 931
          "001111100001" when "011111", -- t[31] = 993
          "010000100001" when "100000", -- t[32] = 1057
          "010001100011" when "100001", -- t[33] = 1123
          "010010100111" when "100010", -- t[34] = 1191
          "010011101101" when "100011", -- t[35] = 1261
          "010100110101" when "100100", -- t[36] = 1333
          "010101111111" when "100101", -- t[37] = 1407
          "010111001011" when "100110", -- t[38] = 1483
          "011000011001" when "100111", -- t[39] = 1561
          "011001101001" when "101000", -- t[40] = 1641
          "011010111010" when "101001", -- t[41] = 1722
          "011100001110" when "101010", -- t[42] = 1806
          "011101100100" when "101011", -- t[43] = 1892
          "011110111100" when "101100", -- t[44] = 1980
          "100000010110" when "101101", -- t[45] = 2070
          "100001110010" when "101110", -- t[46] = 2162
          "100011010000" when "101111", -- t[47] = 2256
          "100100110000" when "110000", -- t[48] = 2352
          "100110010010" when "110001", -- t[49] = 2450
          "100111110111" when "110010", -- t[50] = 2551
          "101001011101" when "110011", -- t[51] = 2653
          "101011000101" when "110100", -- t[52] = 2757
          "101100101111" when "110101", -- t[53] = 2863
          "101110011011" when "110110", -- t[54] = 2971
          "110000001001" when "110111", -- t[55] = 3081
          "110001111001" when "111000", -- t[56] = 3193
          "110011101011" when "111001", -- t[57] = 3307
          "110101011111" when "111010", -- t[58] = 3423
          "110111010101" when "111011", -- t[59] = 3541
          "111001001101" when "111100", -- t[60] = 3661
          "111011000111" when "111101", -- t[61] = 3783
          "111101000011" when "111110", -- t[62] = 3907
          "111111000001" when "111111", -- t[63] = 4033
          "------------" when others;

  r(11 downto 0) <= r0;
  r(12 downto 12) <= (12 downto 12 => ('0'));
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 4; mu_1 = 4; lambda_1 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_21_t1_pow is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_21_t1_pow is
  signal pp0 : std_logic_vector(2 downto 0);
  signal r0 : std_logic_vector(2 downto 0);
begin
  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(2 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 4; sigma'_1,1 = 3; wO_1,1 = 6.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_21_t1_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         s : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_21_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a & s;

  with x select
    r <= "000000" when "0000000", -- t[0] = 0
         "000000" when "0000001", -- t[1] = 0
         "000000" when "0000010", -- t[2] = 0
         "000000" when "0000011", -- t[3] = 0
         "000001" when "0000100", -- t[4] = 1
         "000001" when "0000101", -- t[5] = 1
         "000001" when "0000110", -- t[6] = 1
         "000001" when "0000111", -- t[7] = 1
         "000000" when "0001000", -- t[8] = 0
         "000001" when "0001001", -- t[9] = 1
         "000001" when "0001010", -- t[10] = 1
         "000010" when "0001011", -- t[11] = 2
         "000011" when "0001100", -- t[12] = 3
         "000100" when "0001101", -- t[13] = 4
         "000100" when "0001110", -- t[14] = 4
         "000101" when "0001111", -- t[15] = 5
         "000000" when "0010000", -- t[16] = 0
         "000001" when "0010001", -- t[17] = 1
         "000011" when "0010010", -- t[18] = 3
         "000100" when "0010011", -- t[19] = 4
         "000101" when "0010100", -- t[20] = 5
         "000110" when "0010101", -- t[21] = 6
         "001000" when "0010110", -- t[22] = 8
         "001001" when "0010111", -- t[23] = 9
         "000000" when "0011000", -- t[24] = 0
         "000010" when "0011001", -- t[25] = 2
         "000100" when "0011010", -- t[26] = 4
         "000110" when "0011011", -- t[27] = 6
         "000111" when "0011100", -- t[28] = 7
         "001001" when "0011101", -- t[29] = 9
         "001011" when "0011110", -- t[30] = 11
         "001101" when "0011111", -- t[31] = 13
         "000001" when "0100000", -- t[32] = 1
         "000011" when "0100001", -- t[33] = 3
         "000101" when "0100010", -- t[34] = 5
         "000111" when "0100011", -- t[35] = 7
         "001010" when "0100100", -- t[36] = 10
         "001100" when "0100101", -- t[37] = 12
         "001110" when "0100110", -- t[38] = 14
         "010000" when "0100111", -- t[39] = 16
         "000001" when "0101000", -- t[40] = 1
         "000100" when "0101001", -- t[41] = 4
         "000110" when "0101010", -- t[42] = 6
         "001001" when "0101011", -- t[43] = 9
         "001100" when "0101100", -- t[44] = 12
         "001111" when "0101101", -- t[45] = 15
         "010001" when "0101110", -- t[46] = 17
         "010100" when "0101111", -- t[47] = 20
         "000001" when "0110000", -- t[48] = 1
         "000100" when "0110001", -- t[49] = 4
         "001000" when "0110010", -- t[50] = 8
         "001011" when "0110011", -- t[51] = 11
         "001110" when "0110100", -- t[52] = 14
         "010001" when "0110101", -- t[53] = 17
         "010101" when "0110110", -- t[54] = 21
         "011000" when "0110111", -- t[55] = 24
         "000001" when "0111000", -- t[56] = 1
         "000101" when "0111001", -- t[57] = 5
         "001001" when "0111010", -- t[58] = 9
         "001101" when "0111011", -- t[59] = 13
         "010000" when "0111100", -- t[60] = 16
         "010100" when "0111101", -- t[61] = 20
         "011000" when "0111110", -- t[62] = 24
         "011100" when "0111111", -- t[63] = 28
         "000010" when "1000000", -- t[64] = 2
         "000110" when "1000001", -- t[65] = 6
         "001010" when "1000010", -- t[66] = 10
         "001110" when "1000011", -- t[67] = 14
         "010011" when "1000100", -- t[68] = 19
         "010111" when "1000101", -- t[69] = 23
         "011011" when "1000110", -- t[70] = 27
         "011111" when "1000111", -- t[71] = 31
         "000010" when "1001000", -- t[72] = 2
         "000111" when "1001001", -- t[73] = 7
         "001011" when "1001010", -- t[74] = 11
         "010000" when "1001011", -- t[75] = 16
         "010101" when "1001100", -- t[76] = 21
         "011010" when "1001101", -- t[77] = 26
         "011110" when "1001110", -- t[78] = 30
         "100011" when "1001111", -- t[79] = 35
         "000010" when "1010000", -- t[80] = 2
         "000111" when "1010001", -- t[81] = 7
         "001101" when "1010010", -- t[82] = 13
         "010010" when "1010011", -- t[83] = 18
         "010111" when "1010100", -- t[84] = 23
         "011100" when "1010101", -- t[85] = 28
         "100010" when "1010110", -- t[86] = 34
         "100111" when "1010111", -- t[87] = 39
         "000010" when "1011000", -- t[88] = 2
         "001000" when "1011001", -- t[89] = 8
         "001110" when "1011010", -- t[90] = 14
         "010100" when "1011011", -- t[91] = 20
         "011001" when "1011100", -- t[92] = 25
         "011111" when "1011101", -- t[93] = 31
         "100101" when "1011110", -- t[94] = 37
         "101011" when "1011111", -- t[95] = 43
         "000011" when "1100000", -- t[96] = 3
         "001001" when "1100001", -- t[97] = 9
         "001111" when "1100010", -- t[98] = 15
         "010101" when "1100011", -- t[99] = 21
         "011100" when "1100100", -- t[100] = 28
         "100010" when "1100101", -- t[101] = 34
         "101000" when "1100110", -- t[102] = 40
         "101110" when "1100111", -- t[103] = 46
         "000011" when "1101000", -- t[104] = 3
         "001010" when "1101001", -- t[105] = 10
         "010000" when "1101010", -- t[106] = 16
         "010111" when "1101011", -- t[107] = 23
         "011110" when "1101100", -- t[108] = 30
         "100101" when "1101101", -- t[109] = 37
         "101011" when "1101110", -- t[110] = 43
         "110010" when "1101111", -- t[111] = 50
         "000011" when "1110000", -- t[112] = 3
         "001010" when "1110001", -- t[113] = 10
         "010010" when "1110010", -- t[114] = 18
         "011001" when "1110011", -- t[115] = 25
         "100000" when "1110100", -- t[116] = 32
         "100111" when "1110101", -- t[117] = 39
         "101111" when "1110110", -- t[118] = 47
         "110110" when "1110111", -- t[119] = 54
         "000011" when "1111000", -- t[120] = 3
         "001011" when "1111001", -- t[121] = 11
         "010011" when "1111010", -- t[122] = 19
         "011011" when "1111011", -- t[123] = 27
         "100010" when "1111100", -- t[124] = 34
         "101010" when "1111101", -- t[125] = 42
         "110010" when "1111110", -- t[126] = 50
         "111010" when "1111111", -- t[127] = 58
         "------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 4; beta_1 = 4; lambda_1 = 4;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (ROM):  alpha_1,1 = 4; rho_1,1 = 0; sigma_1,1 = 4; wO_1,1 = 6.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_21_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_21_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(2 downto 0);
  signal s      : std_logic_vector(3 downto 0);
  component fp_exp_exp_y2_21_t1_pow is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  signal a_1    : std_logic_vector(3 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(2 downto 0);
  signal r0_1   : std_logic_vector(5 downto 0);
  signal r_1    : std_logic_vector(12 downto 0);
  component fp_exp_exp_y2_21_t1_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;
begin
  sign <= not b(3);
  b0 <= b(2 downto 0) xor (2 downto 0 => sign);

  pow : fp_exp_exp_y2_21_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(3 downto 0);
  sign_1 <= not s(3);
  s_1 <= s(2 downto 0) xor (2 downto 0 => sign_1);
  t_1 : fp_exp_exp_y2_21_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_1 );
  r_1(5 downto 0) <=
    r0_1 xor (5 downto 0 => ((sign xor sign_1)));
  r_1(12 downto 6) <= (12 downto 6 => ((sign xor sign_1)));

  r <= r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_21_t1_clk is
  port ( a   : in  std_logic_vector(3 downto 0);
         b   : in  std_logic_vector(3 downto 0);
         r   : out std_logic_vector(12 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_21_t1_clk is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(2 downto 0);
  signal s      : std_logic_vector(3 downto 0);
  component fp_exp_exp_y2_21_t1_pow is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  signal a_1     : std_logic_vector(3 downto 0);
  signal sign_1  : std_logic;
  signal s_1     : std_logic_vector(2 downto 0);
  signal r0_10   : std_logic_vector(5 downto 0);
  signal r0_1r   : std_logic_vector(5 downto 0);
  signal r_1     : std_logic_vector(12 downto 0);
  signal sign_10 : std_logic;
  signal sign_1r : std_logic;
  component fp_exp_exp_y2_21_t1_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;
begin
  sign <= not b(3);
  b0 <= b(2 downto 0) xor (2 downto 0 => sign);

  pow : fp_exp_exp_y2_21_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(3 downto 0);
  sign_1 <= not s(3);
  s_1 <= s(2 downto 0) xor (2 downto 0 => sign_1);
  sign_10 <= sign xor sign_1;
  t_1 : fp_exp_exp_y2_21_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_10 );
  r_1(5 downto 0) <=
    r0_1r xor (5 downto 0 => sign_1r);
  r_1(12 downto 6) <= (12 downto 6 => sign_1r);

  process(clk)
  begin
    if clk'event and clk = '1' then
      r0_1r   <= r0_10;
      sign_1r <= sign_10;
    end if;
  end process;

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_21 is
  port ( x : in  std_logic_vector(9 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_21 is
  signal a_0 : std_logic_vector(5 downto 0);
  signal r_0 : std_logic_vector(12 downto 0);
  component fp_exp_exp_y2_21_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  signal a_1 : std_logic_vector(3 downto 0);
  signal b_1 : std_logic_vector(3 downto 0);
  signal r_1 : std_logic_vector(12 downto 0);
  component fp_exp_exp_y2_21_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  signal sum : std_logic_vector(12 downto 0);
begin
  a_0 <= x(9 downto 4);
  t_0 : fp_exp_exp_y2_21_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(9 downto 6);
  b_1 <= x(3 downto 0);
  t_1 : fp_exp_exp_y2_21_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  sum <= r_0 + r_1;
  r <= sum(12 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_21_clk is
  port ( x   : in  std_logic_vector(9 downto 0);
         r   : out std_logic_vector(10 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_21_clk is
  signal a_x0 : std_logic_vector(5 downto 0);
  signal a_xr : std_logic_vector(5 downto 0);
  signal r_0  : std_logic_vector(12 downto 0);
  component fp_exp_exp_y2_21_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  signal a_1 : std_logic_vector(3 downto 0);
  signal b_1 : std_logic_vector(3 downto 0);
  signal r_1 : std_logic_vector(12 downto 0);
  component fp_exp_exp_y2_21_t1_clk is
    port ( a   : in  std_logic_vector(3 downto 0);
           b   : in  std_logic_vector(3 downto 0);
           r   : out std_logic_vector(12 downto 0);
           clk : in  std_logic );
  end component;

  signal sum : std_logic_vector(12 downto 0);
begin
  a_x0 <= x(9 downto 4);
  t_0 : fp_exp_exp_y2_21_t0
    port map ( a => a_xr,
               r => r_0 );

  process(clk)
  begin
    if clk'event and clk = '1' then
      a_xr <= a_x0;
    end if;
  end process;

  a_1 <= x(9 downto 6);
  b_1 <= x(3 downto 0);
  t_1 : fp_exp_exp_y2_21_t1_clk
    port map ( a   => a_1,
               b   => b_1,
               r   => r_1,
               clk => clk );

  sum <= r_0 + r_1;
  r <= sum(12 downto 2);
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function e^x-x-1.
-- wI = 11; wO = 11.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 6; beta = 5;
--   T_0 (ROM):     alpha_0 = 6; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 5; beta_1 = 5.
-- Guard bits: g = 2.
-- Command line: exp 11 11 1   rom 6 0   pm 5 5  ah 5 5 5  0 2  5 3 0  3 2 3


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 6; beta_0 = 0; wO_0 = 13.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22_t0 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_22_t0 is
  signal x0   : std_logic_vector(5 downto 0);
  signal r0   : std_logic_vector(12 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "0000000000011" when "000000", -- t[0] = 3
          "0000000000111" when "000001", -- t[1] = 7
          "0000000001111" when "000010", -- t[2] = 15
          "0000000011011" when "000011", -- t[3] = 27
          "0000000101011" when "000100", -- t[4] = 43
          "0000000111111" when "000101", -- t[5] = 63
          "0000001010111" when "000110", -- t[6] = 87
          "0000001110011" when "000111", -- t[7] = 115
          "0000010010011" when "001000", -- t[8] = 147
          "0000010110111" when "001001", -- t[9] = 183
          "0000011011111" when "001010", -- t[10] = 223
          "0000100001011" when "001011", -- t[11] = 267
          "0000100111010" when "001100", -- t[12] = 314
          "0000101101110" when "001101", -- t[13] = 366
          "0000110100110" when "001110", -- t[14] = 422
          "0000111100010" when "001111", -- t[15] = 482
          "0001000100010" when "010000", -- t[16] = 546
          "0001001100110" when "010001", -- t[17] = 614
          "0001010101110" when "010010", -- t[18] = 686
          "0001011111010" when "010011", -- t[19] = 762
          "0001101001010" when "010100", -- t[20] = 842
          "0001110011110" when "010101", -- t[21] = 926
          "0001111110110" when "010110", -- t[22] = 1014
          "0010001010010" when "010111", -- t[23] = 1106
          "0010010110010" when "011000", -- t[24] = 1202
          "0010100010110" when "011001", -- t[25] = 1302
          "0010101111110" when "011010", -- t[26] = 1406
          "0010111101010" when "011011", -- t[27] = 1514
          "0011001011010" when "011100", -- t[28] = 1626
          "0011011001110" when "011101", -- t[29] = 1742
          "0011101000110" when "011110", -- t[30] = 1862
          "0011111000010" when "011111", -- t[31] = 1986
          "0100001000010" when "100000", -- t[32] = 2114
          "0100011000110" when "100001", -- t[33] = 2246
          "0100101001110" when "100010", -- t[34] = 2382
          "0100111011010" when "100011", -- t[35] = 2522
          "0101001101010" when "100100", -- t[36] = 2666
          "0101011111110" when "100101", -- t[37] = 2814
          "0101110010110" when "100110", -- t[38] = 2966
          "0110000110010" when "100111", -- t[39] = 3122
          "0110011010010" when "101000", -- t[40] = 3282
          "0110101110110" when "101001", -- t[41] = 3446
          "0111000011110" when "101010", -- t[42] = 3614
          "0111011001010" when "101011", -- t[43] = 3786
          "0111101111010" when "101100", -- t[44] = 3962
          "1000000101110" when "101101", -- t[45] = 4142
          "1000011100110" when "101110", -- t[46] = 4326
          "1000110100010" when "101111", -- t[47] = 4514
          "1001001100011" when "110000", -- t[48] = 4707
          "1001100100111" when "110001", -- t[49] = 4903
          "1001111101111" when "110010", -- t[50] = 5103
          "1010010111011" when "110011", -- t[51] = 5307
          "1010110001011" when "110100", -- t[52] = 5515
          "1011001011111" when "110101", -- t[53] = 5727
          "1011100110111" when "110110", -- t[54] = 5943
          "1100000010011" when "110111", -- t[55] = 6163
          "1100011110011" when "111000", -- t[56] = 6387
          "1100111011000" when "111001", -- t[57] = 6616
          "1101011000000" when "111010", -- t[58] = 6848
          "1101110101100" when "111011", -- t[59] = 7084
          "1110010011100" when "111100", -- t[60] = 7324
          "1110110010000" when "111101", -- t[61] = 7568
          "1111010001000" when "111110", -- t[62] = 7816
          "1111110000100" when "111111", -- t[63] = 8068
          "-------------" when others;

  r(12 downto 0) <= r0;
  r(13 downto 13) <= (13 downto 13 => ('0'));
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 5; mu_1 = 5; lambda_1 = 5.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22_t1_pow is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_22_t1_pow is
  signal pp0 : std_logic_vector(3 downto 0);
  signal r0 : std_logic_vector(3 downto 0);
begin
  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(3 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 5; sigma'_1,1 = 2; wO_1,1 = 7.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22_t1_t1 is
  port ( a : in  std_logic_vector(4 downto 0);
         s : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_22_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0000000" when "0000000", -- t[0] = 0
         "0000000" when "0000001", -- t[1] = 0
         "0000001" when "0000010", -- t[2] = 1
         "0000001" when "0000011", -- t[3] = 1
         "0000000" when "0000100", -- t[4] = 0
         "0000010" when "0000101", -- t[5] = 2
         "0000011" when "0000110", -- t[6] = 3
         "0000101" when "0000111", -- t[7] = 5
         "0000001" when "0001000", -- t[8] = 1
         "0000011" when "0001001", -- t[9] = 3
         "0000110" when "0001010", -- t[10] = 6
         "0001000" when "0001011", -- t[11] = 8
         "0000001" when "0001100", -- t[12] = 1
         "0000101" when "0001101", -- t[13] = 5
         "0001000" when "0001110", -- t[14] = 8
         "0001100" when "0001111", -- t[15] = 12
         "0000010" when "0010000", -- t[16] = 2
         "0000110" when "0010001", -- t[17] = 6
         "0001011" when "0010010", -- t[18] = 11
         "0001111" when "0010011", -- t[19] = 15
         "0000010" when "0010100", -- t[20] = 2
         "0001000" when "0010101", -- t[21] = 8
         "0001101" when "0010110", -- t[22] = 13
         "0010011" when "0010111", -- t[23] = 19
         "0000011" when "0011000", -- t[24] = 3
         "0001001" when "0011001", -- t[25] = 9
         "0010000" when "0011010", -- t[26] = 16
         "0010110" when "0011011", -- t[27] = 22
         "0000011" when "0011100", -- t[28] = 3
         "0001011" when "0011101", -- t[29] = 11
         "0010010" when "0011110", -- t[30] = 18
         "0011010" when "0011111", -- t[31] = 26
         "0000100" when "0100000", -- t[32] = 4
         "0001100" when "0100001", -- t[33] = 12
         "0010101" when "0100010", -- t[34] = 21
         "0011101" when "0100011", -- t[35] = 29
         "0000100" when "0100100", -- t[36] = 4
         "0001110" when "0100101", -- t[37] = 14
         "0010111" when "0100110", -- t[38] = 23
         "0100001" when "0100111", -- t[39] = 33
         "0000101" when "0101000", -- t[40] = 5
         "0001111" when "0101001", -- t[41] = 15
         "0011010" when "0101010", -- t[42] = 26
         "0100100" when "0101011", -- t[43] = 36
         "0000101" when "0101100", -- t[44] = 5
         "0010001" when "0101101", -- t[45] = 17
         "0011100" when "0101110", -- t[46] = 28
         "0101000" when "0101111", -- t[47] = 40
         "0000110" when "0110000", -- t[48] = 6
         "0010010" when "0110001", -- t[49] = 18
         "0011111" when "0110010", -- t[50] = 31
         "0101011" when "0110011", -- t[51] = 43
         "0000110" when "0110100", -- t[52] = 6
         "0010100" when "0110101", -- t[53] = 20
         "0100001" when "0110110", -- t[54] = 33
         "0101111" when "0110111", -- t[55] = 47
         "0000111" when "0111000", -- t[56] = 7
         "0010101" when "0111001", -- t[57] = 21
         "0100100" when "0111010", -- t[58] = 36
         "0110010" when "0111011", -- t[59] = 50
         "0000111" when "0111100", -- t[60] = 7
         "0010111" when "0111101", -- t[61] = 23
         "0100110" when "0111110", -- t[62] = 38
         "0110110" when "0111111", -- t[63] = 54
         "0001000" when "1000000", -- t[64] = 8
         "0011000" when "1000001", -- t[65] = 24
         "0101001" when "1000010", -- t[66] = 41
         "0111001" when "1000011", -- t[67] = 57
         "0001000" when "1000100", -- t[68] = 8
         "0011010" when "1000101", -- t[69] = 26
         "0101011" when "1000110", -- t[70] = 43
         "0111101" when "1000111", -- t[71] = 61
         "0001001" when "1001000", -- t[72] = 9
         "0011011" when "1001001", -- t[73] = 27
         "0101110" when "1001010", -- t[74] = 46
         "1000000" when "1001011", -- t[75] = 64
         "0001001" when "1001100", -- t[76] = 9
         "0011101" when "1001101", -- t[77] = 29
         "0110000" when "1001110", -- t[78] = 48
         "1000100" when "1001111", -- t[79] = 68
         "0001010" when "1010000", -- t[80] = 10
         "0011110" when "1010001", -- t[81] = 30
         "0110011" when "1010010", -- t[82] = 51
         "1000111" when "1010011", -- t[83] = 71
         "0001010" when "1010100", -- t[84] = 10
         "0100000" when "1010101", -- t[85] = 32
         "0110101" when "1010110", -- t[86] = 53
         "1001011" when "1010111", -- t[87] = 75
         "0001011" when "1011000", -- t[88] = 11
         "0100001" when "1011001", -- t[89] = 33
         "0111000" when "1011010", -- t[90] = 56
         "1001110" when "1011011", -- t[91] = 78
         "0001011" when "1011100", -- t[92] = 11
         "0100011" when "1011101", -- t[93] = 35
         "0111010" when "1011110", -- t[94] = 58
         "1010010" when "1011111", -- t[95] = 82
         "0001100" when "1100000", -- t[96] = 12
         "0100100" when "1100001", -- t[97] = 36
         "0111101" when "1100010", -- t[98] = 61
         "1010101" when "1100011", -- t[99] = 85
         "0001100" when "1100100", -- t[100] = 12
         "0100110" when "1100101", -- t[101] = 38
         "0111111" when "1100110", -- t[102] = 63
         "1011001" when "1100111", -- t[103] = 89
         "0001101" when "1101000", -- t[104] = 13
         "0100111" when "1101001", -- t[105] = 39
         "1000010" when "1101010", -- t[106] = 66
         "1011100" when "1101011", -- t[107] = 92
         "0001101" when "1101100", -- t[108] = 13
         "0101001" when "1101101", -- t[109] = 41
         "1000100" when "1101110", -- t[110] = 68
         "1100000" when "1101111", -- t[111] = 96
         "0001110" when "1110000", -- t[112] = 14
         "0101010" when "1110001", -- t[113] = 42
         "1000111" when "1110010", -- t[114] = 71
         "1100011" when "1110011", -- t[115] = 99
         "0001110" when "1110100", -- t[116] = 14
         "0101100" when "1110101", -- t[117] = 44
         "1001001" when "1110110", -- t[118] = 73
         "1100111" when "1110111", -- t[119] = 103
         "0001111" when "1111000", -- t[120] = 15
         "0101101" when "1111001", -- t[121] = 45
         "1001100" when "1111010", -- t[122] = 76
         "1101010" when "1111011", -- t[123] = 106
         "0001111" when "1111100", -- t[124] = 15
         "0101111" when "1111101", -- t[125] = 47
         "1001110" when "1111110", -- t[126] = 78
         "1101110" when "1111111", -- t[127] = 110
         "-------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_2.
-- Decomposition:
--   alpha_1,2 = 3; sigma'_1,2 = 1; wO_1,2 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22_t1_t2 is
  port ( a : in  std_logic_vector(2 downto 0);
         s : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_22_t1_t2 is
  signal x : std_logic_vector(3 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0000" when "0000", -- t[0] = 0
         "0000" when "0001", -- t[1] = 0
         "0000" when "0010", -- t[2] = 0
         "0010" when "0011", -- t[3] = 2
         "0001" when "0100", -- t[4] = 1
         "0011" when "0101", -- t[5] = 3
         "0001" when "0110", -- t[6] = 1
         "0101" when "0111", -- t[7] = 5
         "0010" when "1000", -- t[8] = 2
         "0110" when "1001", -- t[9] = 6
         "0010" when "1010", -- t[10] = 2
         "1000" when "1011", -- t[11] = 8
         "0011" when "1100", -- t[12] = 3
         "1001" when "1101", -- t[13] = 9
         "0011" when "1110", -- t[14] = 3
         "1011" when "1111", -- t[15] = 11
         "----" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 5; beta_1 = 5; lambda_1 = 5;  m_1 = 2;
--   Pow   (AdHoc);
--   Q_1,1 (ROM):  alpha_1,1 = 5; rho_1,1 = 0; sigma_1,1 = 3; wO_1,1 = 7;
--   Q_1,2 (ROM):  alpha_1,2 = 3; rho_1,2 = 3; sigma_1,2 = 2; wO_1,2 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22_t1 is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_22_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(3 downto 0);
  signal s      : std_logic_vector(4 downto 0);
  component fp_exp_exp_y2_22_t1_pow is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;

  signal a_1    : std_logic_vector(4 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(1 downto 0);
  signal r0_1   : std_logic_vector(6 downto 0);
  signal r_1    : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_22_t1_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           s : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  signal a_2    : std_logic_vector(2 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(0 downto 0);
  signal r0_2   : std_logic_vector(3 downto 0);
  signal r_2    : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_22_t1_t2 is
    port ( a : in  std_logic_vector(2 downto 0);
           s : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;
begin
  sign <= not b(4);
  b0 <= b(3 downto 0) xor (3 downto 0 => sign);

  pow : fp_exp_exp_y2_22_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(4 downto 0);
  sign_1 <= not s(4);
  s_1 <= s(3 downto 2) xor (3 downto 2 => sign_1);
  t_1 : fp_exp_exp_y2_22_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_1 );
  r_1(6 downto 0) <=
    r0_1 xor (6 downto 0 => ((sign xor sign_1)));
  r_1(13 downto 7) <= (13 downto 7 => ((sign xor sign_1)));

  a_2 <= a(4 downto 2);
  sign_2 <= not s(1);
  s_2 <= s(0 downto 0) xor (0 downto 0 => sign_2);
  t_2 : fp_exp_exp_y2_22_t1_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(3 downto 0) <=
    r0_2 xor (3 downto 0 => ((sign xor sign_2)));
  r_2(13 downto 4) <= (13 downto 4 => ((sign xor sign_2)));

  r <= r_1 + r_2;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22_t1_clk is
  port ( a   : in  std_logic_vector(4 downto 0);
         b   : in  std_logic_vector(4 downto 0);
         r   : out std_logic_vector(13 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_22_t1_clk is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(3 downto 0);
  signal s      : std_logic_vector(4 downto 0);
  component fp_exp_exp_y2_22_t1_pow is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;

  signal a_1     : std_logic_vector(4 downto 0);
  signal sign_1  : std_logic;
  signal s_1     : std_logic_vector(1 downto 0);
  signal r0_10   : std_logic_vector(6 downto 0);
  signal r0_1r   : std_logic_vector(6 downto 0);
  signal r_1     : std_logic_vector(13 downto 0);
  signal sign_10 : std_logic;
  signal sign_1r : std_logic;
  component fp_exp_exp_y2_22_t1_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           s : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  signal a_2     : std_logic_vector(2 downto 0);
  signal sign_2  : std_logic;
  signal s_2     : std_logic_vector(0 downto 0);
  signal r0_20   : std_logic_vector(3 downto 0);
  signal r0_2r   : std_logic_vector(3 downto 0);
  signal r_2     : std_logic_vector(13 downto 0);
  signal sign_20 : std_logic;
  signal sign_2r : std_logic;
  component fp_exp_exp_y2_22_t1_t2 is
    port ( a : in  std_logic_vector(2 downto 0);
           s : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;
begin
  sign <= not b(4);
  b0 <= b(3 downto 0) xor (3 downto 0 => sign);

  pow : fp_exp_exp_y2_22_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(4 downto 0);
  sign_1 <= not s(4);
  s_1 <= s(3 downto 2) xor (3 downto 2 => sign_1);
  sign_10 <= sign xor sign_1;
  t_1 : fp_exp_exp_y2_22_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_10 );
  r_1(6 downto 0) <=
    r0_1r xor (6 downto 0 => sign_1r);
  r_1(13 downto 7) <= (13 downto 7 => sign_1r);

  a_2 <= a(4 downto 2);
  sign_2 <= not s(1);
  s_2 <= s(0 downto 0) xor (0 downto 0 => sign_2);
  sign_20 <= sign xor sign_2;
  t_2 : fp_exp_exp_y2_22_t1_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_20 );
  r_2(3 downto 0) <=
    r0_2r xor (3 downto 0 => sign_2r);
  r_2(13 downto 4) <= (13 downto 4 => sign_2r);

  process(clk)
  begin
    if clk'event and clk = '1' then
      r0_1r   <= r0_10;
      sign_1r <= sign_10;
      r0_2r   <= r0_20;
      sign_2r <= sign_20;
    end if;
  end process;
  
  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22 is
  port ( x : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_22 is
  signal a_0 : std_logic_vector(5 downto 0);
  signal r_0 : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_22_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1 : std_logic_vector(4 downto 0);
  signal b_1 : std_logic_vector(4 downto 0);
  signal r_1 : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_22_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal sum : std_logic_vector(13 downto 0);
begin
  a_0 <= x(10 downto 5);
  t_0 : fp_exp_exp_y2_22_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(10 downto 6);
  b_1 <= x(4 downto 0);
  t_1 : fp_exp_exp_y2_22_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  sum <= r_0 + r_1;
  r <= sum(13 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_22_clk is
  port ( x   : in  std_logic_vector(10 downto 0);
         r   : out std_logic_vector(11 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_22_clk is
  signal a_x0 : std_logic_vector(5 downto 0);
  signal a_xr : std_logic_vector(5 downto 0);
  signal r_0  : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_22_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1 : std_logic_vector(4 downto 0);
  signal b_1 : std_logic_vector(4 downto 0);
  signal r_1 : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_22_t1_clk is
    port ( a   : in  std_logic_vector(4 downto 0);
           b   : in  std_logic_vector(4 downto 0);
           r   : out std_logic_vector(13 downto 0);
           clk : in  std_logic );
  end component;

  signal sum : std_logic_vector(13 downto 0);
begin
  a_x0 <= x(10 downto 5);
  t_0 : fp_exp_exp_y2_22_t0
    port map ( a => a_xr,
               r => r_0 );

  process(clk)
  begin
    if clk'event and clk = '1' then
      a_xr <= a_x0;
    end if;
  end process;

  a_1 <= x(10 downto 6);
  b_1 <= x(4 downto 0);
  t_1 : fp_exp_exp_y2_22_t1_clk
    port map ( a   => a_1,
               b   => b_1,
               r   => r_1,
               clk => clk );

  sum <= r_0 + r_1;
  r <= sum(13 downto 2);
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function e^x-x-1.
-- wI = 12; wO = 12.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 6; beta = 6;
--   T_0 (ROM):     alpha_0 = 6; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 6; beta_1 = 6.
-- Guard bits: g = 1.
-- Command line: exp 12 12 1   rom 6 0   pm 6 6  ah 6 6 6  1 0  6 6 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 6; beta_0 = 0; wO_0 = 13.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_23_t0 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_23_t0 is
  signal x0   : std_logic_vector(5 downto 0);
  signal r0   : std_logic_vector(12 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "0000000000010" when "000000", -- t[0] = 2
          "0000000000110" when "000001", -- t[1] = 6
          "0000000001110" when "000010", -- t[2] = 14
          "0000000011010" when "000011", -- t[3] = 26
          "0000000101010" when "000100", -- t[4] = 42
          "0000000111110" when "000101", -- t[5] = 62
          "0000001010110" when "000110", -- t[6] = 86
          "0000001110010" when "000111", -- t[7] = 114
          "0000010010001" when "001000", -- t[8] = 145
          "0000010110101" when "001001", -- t[9] = 181
          "0000011011101" when "001010", -- t[10] = 221
          "0000100001001" when "001011", -- t[11] = 265
          "0000100111001" when "001100", -- t[12] = 313
          "0000101101101" when "001101", -- t[13] = 365
          "0000110100101" when "001110", -- t[14] = 421
          "0000111100001" when "001111", -- t[15] = 481
          "0001000100001" when "010000", -- t[16] = 545
          "0001001100101" when "010001", -- t[17] = 613
          "0001010101101" when "010010", -- t[18] = 685
          "0001011111001" when "010011", -- t[19] = 761
          "0001101001001" when "010100", -- t[20] = 841
          "0001110011101" when "010101", -- t[21] = 925
          "0001111110101" when "010110", -- t[22] = 1013
          "0010001010001" when "010111", -- t[23] = 1105
          "0010010110001" when "011000", -- t[24] = 1201
          "0010100010101" when "011001", -- t[25] = 1301
          "0010101111101" when "011010", -- t[26] = 1405
          "0010111101001" when "011011", -- t[27] = 1513
          "0011001011001" when "011100", -- t[28] = 1625
          "0011011001101" when "011101", -- t[29] = 1741
          "0011101000101" when "011110", -- t[30] = 1861
          "0011111000001" when "011111", -- t[31] = 1985
          "0100001000001" when "100000", -- t[32] = 2113
          "0100011000101" when "100001", -- t[33] = 2245
          "0100101001101" when "100010", -- t[34] = 2381
          "0100111011010" when "100011", -- t[35] = 2522
          "0101001101010" when "100100", -- t[36] = 2666
          "0101011111110" when "100101", -- t[37] = 2814
          "0101110010110" when "100110", -- t[38] = 2966
          "0110000110010" when "100111", -- t[39] = 3122
          "0110011010010" when "101000", -- t[40] = 3282
          "0110101110110" when "101001", -- t[41] = 3446
          "0111000011110" when "101010", -- t[42] = 3614
          "0111011001010" when "101011", -- t[43] = 3786
          "0111101111010" when "101100", -- t[44] = 3962
          "1000000101110" when "101101", -- t[45] = 4142
          "1000011100110" when "101110", -- t[46] = 4326
          "1000110100010" when "101111", -- t[47] = 4514
          "1001001100011" when "110000", -- t[48] = 4707
          "1001100100111" when "110001", -- t[49] = 4903
          "1001111101111" when "110010", -- t[50] = 5103
          "1010010111011" when "110011", -- t[51] = 5307
          "1010110001011" when "110100", -- t[52] = 5515
          "1011001011111" when "110101", -- t[53] = 5727
          "1011100110111" when "110110", -- t[54] = 5943
          "1100000010011" when "110111", -- t[55] = 6163
          "1100011110100" when "111000", -- t[56] = 6388
          "1100111011000" when "111001", -- t[57] = 6616
          "1101011000000" when "111010", -- t[58] = 6848
          "1101110101100" when "111011", -- t[59] = 7084
          "1110010011100" when "111100", -- t[60] = 7324
          "1110110010001" when "111101", -- t[61] = 7569
          "1111010001001" when "111110", -- t[62] = 7817
          "1111110000101" when "111111", -- t[63] = 8069
          "-------------" when others;

  r(12 downto 0) <= r0;
  r(13 downto 13) <= (13 downto 13 => ('0'));
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 6; mu_1 = 6; lambda_1 = 6.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_23_t1_pow is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_23_t1_pow is
  signal pp0 : std_logic_vector(4 downto 0);
  signal r0 : std_logic_vector(4 downto 0);
begin
  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(4 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 6; wO_1,1 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_23_t1_t1 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_23_t1_t1 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a;

  with x select
    r <= "00000010" when "000000", -- t[0] = 2
         "00000110" when "000001", -- t[1] = 6
         "00001010" when "000010", -- t[2] = 10
         "00001110" when "000011", -- t[3] = 14
         "00010010" when "000100", -- t[4] = 18
         "00010110" when "000101", -- t[5] = 22
         "00011010" when "000110", -- t[6] = 26
         "00011110" when "000111", -- t[7] = 30
         "00100010" when "001000", -- t[8] = 34
         "00100110" when "001001", -- t[9] = 38
         "00101010" when "001010", -- t[10] = 42
         "00101110" when "001011", -- t[11] = 46
         "00110010" when "001100", -- t[12] = 50
         "00110110" when "001101", -- t[13] = 54
         "00111010" when "001110", -- t[14] = 58
         "00111110" when "001111", -- t[15] = 62
         "01000010" when "010000", -- t[16] = 66
         "01000110" when "010001", -- t[17] = 70
         "01001010" when "010010", -- t[18] = 74
         "01001110" when "010011", -- t[19] = 78
         "01010010" when "010100", -- t[20] = 82
         "01010110" when "010101", -- t[21] = 86
         "01011010" when "010110", -- t[22] = 90
         "01011110" when "010111", -- t[23] = 94
         "01100010" when "011000", -- t[24] = 98
         "01100110" when "011001", -- t[25] = 102
         "01101010" when "011010", -- t[26] = 106
         "01101110" when "011011", -- t[27] = 110
         "01110010" when "011100", -- t[28] = 114
         "01110110" when "011101", -- t[29] = 118
         "01111010" when "011110", -- t[30] = 122
         "01111110" when "011111", -- t[31] = 126
         "10000010" when "100000", -- t[32] = 130
         "10000110" when "100001", -- t[33] = 134
         "10001010" when "100010", -- t[34] = 138
         "10001110" when "100011", -- t[35] = 142
         "10010010" when "100100", -- t[36] = 146
         "10010110" when "100101", -- t[37] = 150
         "10011010" when "100110", -- t[38] = 154
         "10011110" when "100111", -- t[39] = 158
         "10100010" when "101000", -- t[40] = 162
         "10100110" when "101001", -- t[41] = 166
         "10101010" when "101010", -- t[42] = 170
         "10101110" when "101011", -- t[43] = 174
         "10110010" when "101100", -- t[44] = 178
         "10110110" when "101101", -- t[45] = 182
         "10111010" when "101110", -- t[46] = 186
         "10111110" when "101111", -- t[47] = 190
         "11000010" when "110000", -- t[48] = 194
         "11000110" when "110001", -- t[49] = 198
         "11001010" when "110010", -- t[50] = 202
         "11001110" when "110011", -- t[51] = 206
         "11010010" when "110100", -- t[52] = 210
         "11010110" when "110101", -- t[53] = 214
         "11011010" when "110110", -- t[54] = 218
         "11011110" when "110111", -- t[55] = 222
         "11100010" when "111000", -- t[56] = 226
         "11100110" when "111001", -- t[57] = 230
         "11101010" when "111010", -- t[58] = 234
         "11101110" when "111011", -- t[59] = 238
         "11110010" when "111100", -- t[60] = 242
         "11110110" when "111101", -- t[61] = 246
         "11111010" when "111110", -- t[62] = 250
         "11111110" when "111111", -- t[63] = 254
         "--------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 6; beta_1 = 6; lambda_1 = 6;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 6; rho_1,1 = 0; sigma_1,1 = 6; wO_1,1 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_23_t1 is
  port ( a : in  std_logic_vector(5 downto 0);
         b : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_23_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(4 downto 0);
  signal s      : std_logic_vector(5 downto 0);
  component fp_exp_exp_y2_23_t1_pow is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  signal a_1    : std_logic_vector(5 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(4 downto 0);
  signal k_1    : std_logic_vector(7 downto 0);
  signal r0_1   : std_logic_vector(14 downto 0);
  signal r_1    : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_23_t1_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;
begin
  sign <= not b(5);
  b0 <= b(4 downto 0) xor (4 downto 0 => sign);

  pow : fp_exp_exp_y2_23_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(5 downto 0);
  sign_1 <= not s(5);
  s_1 <= s(4 downto 0) xor (4 downto 0 => sign_1);
  t_1 : fp_exp_exp_y2_23_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(7 downto 0) <=
    r0_1(14 downto 7) xor (14 downto 7 => ((sign xor sign_1)));
  r_1(13 downto 8) <= (13 downto 8 => ((sign xor sign_1)));

  r <= r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library work;
use work.pkg_fp_exp.all;

entity fp_exp_exp_y2_23_t1_clk is
  port ( a   : in  std_logic_vector(5 downto 0);
         b   : in  std_logic_vector(5 downto 0);
         r   : out std_logic_vector(13 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_23_t1_clk is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(4 downto 0);
  signal s      : std_logic_vector(5 downto 0);
  component fp_exp_exp_y2_23_t1_pow is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  signal a_1     : std_logic_vector(5 downto 0);
  signal sign_1  : std_logic;
  signal s_1     : std_logic_vector(5 downto 0);
  signal k_1     : std_logic_vector(7 downto 0);
  signal r0_1    : std_logic_vector(14 downto 0);
  signal r_1     : std_logic_vector(13 downto 0);
  signal sign_x0 : std_logic;
  signal sign_xr : std_logic;
  component fp_exp_exp_y2_23_t1_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;
begin
  sign <= not b(5);
  b0 <= b(4 downto 0) xor (4 downto 0 => sign);

  pow : fp_exp_exp_y2_23_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(5 downto 0);
  sign_1 <= not s(5);
  s_1 <= "1" & (s(4 downto 0) xor (4 downto 0 => sign_1));
  t_1 : fp_exp_exp_y2_23_t1_t1
    port map ( a => a_1,
               r => k_1 );

  mult_r0_1 : mult_clk
    generic map ( wX    => 8,
                  wY    => 6,
                  first => 1,
                  steps => 3 )
    port map ( nX  => k_1,
               nY  => s_1,
               nR  => r0_1(13 downto 0),
               clk => clk );
  r0_1(14) <= '0';

  sign_x0 <= sign xor sign_1;
  process(clk)
  begin
    if clk'event and clk = '1' then
      sign_xr <= sign_x0;
    end if;
  end process;

  r_1(7 downto 0) <=
    r0_1(14 downto 7) xor (14 downto 7 => sign_xr);
  r_1(13 downto 8) <= (13 downto 8 => sign_xr);

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_23 is
  port ( x : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of fp_exp_exp_y2_23 is
  signal a_0 : std_logic_vector(5 downto 0);
  signal r_0 : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_23_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1 : std_logic_vector(5 downto 0);
  signal b_1 : std_logic_vector(5 downto 0);
  signal r_1 : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_23_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           b : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal sum : std_logic_vector(13 downto 0);
begin
  a_0 <= x(11 downto 6);
  t_0 : fp_exp_exp_y2_23_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(11 downto 6);
  b_1 <= x(5 downto 0);
  t_1 : fp_exp_exp_y2_23_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  sum <= r_0 + r_1;
  r <= sum(13 downto 1);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_exp_exp_y2_23_clk is
  port ( x   : in  std_logic_vector(11 downto 0);
         r   : out std_logic_vector(12 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_23_clk is
  signal a_x0 : std_logic_vector(5 downto 0);
  signal a_xr : std_logic_vector(5 downto 0);
  signal r_0  : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_23_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1 : std_logic_vector(5 downto 0);
  signal b_1 : std_logic_vector(5 downto 0);
  signal r_1 : std_logic_vector(13 downto 0);
  component fp_exp_exp_y2_23_t1_clk is
    port ( a   : in  std_logic_vector(5 downto 0);
           b   : in  std_logic_vector(5 downto 0);
           r   : out std_logic_vector(13 downto 0);
           clk : in  std_logic );
  end component;

  signal sum : std_logic_vector(13 downto 0);
begin
  a_x0 <= x(11 downto 6);
  t_0 : fp_exp_exp_y2_23_t0
    port map ( a => a_xr,
               r => r_0 );

  process(clk)
  begin
    if clk'event and clk = '1' then
      a_xr <= a_x0;
    end if;
  end process;

  a_1 <= x(11 downto 6);
  b_1 <= x(5 downto 0);
  t_1 : fp_exp_exp_y2_23_t1_clk
    port map ( a   => a_1,
               b   => b_1,
               r   => r_1,
               clk => clk );

  sum <= r_0 + r_1;
  r <= sum(13 downto 1);
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library work;
use work.pkg_fp_exp.all;
use work.pkg_fp_exp_exp_y2.all;

entity fp_exp_exp_y2 is
  generic ( wF : positive );
  port ( nY2    : in  std_logic_vector(fp_exp_wy2(wF)-1 downto 0);
         nExpY2 : out std_logic_vector(fp_exp_wy2(wF) downto 0) );
end entity;

architecture arch of fp_exp_exp_y2 is
begin

  exp_y2_6 : if wF = 6 generate
    exp_y2 : fp_exp_exp_y2_6
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_7 : if wF = 7 generate
    exp_y2 : fp_exp_exp_y2_7
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_8 : if wF = 8 generate
    exp_y2 : fp_exp_exp_y2_8
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_9 : if wF = 9 generate
    exp_y2 : fp_exp_exp_y2_9
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_10 : if wF = 10 generate
    exp_y2 : fp_exp_exp_y2_10
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_11 : if wF = 11 generate
    exp_y2 : fp_exp_exp_y2_11
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_12 : if wF = 12 generate
    exp_y2 : fp_exp_exp_y2_12
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_13 : if wF = 13 generate
    exp_y2 : fp_exp_exp_y2_13
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_14 : if wF = 14 generate
    exp_y2 : fp_exp_exp_y2_14
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_15 : if wF = 15 generate
    exp_y2 : fp_exp_exp_y2_15
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_16 : if wF = 16 generate
    exp_y2 : fp_exp_exp_y2_16
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_17 : if wF = 17 generate
    exp_y2 : fp_exp_exp_y2_17
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_18 : if wF = 18 generate
    exp_y2 : fp_exp_exp_y2_18
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_19 : if wF = 19 generate
    exp_y2 : fp_exp_exp_y2_19
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_20 : if wF = 20 generate
    exp_y2 : fp_exp_exp_y2_20
      port map ( x => nY2,
                 r => nExpY2 );
  end generate;

  exp_y2_21 : if wF = 21 generate
    exp_y2 : fp_exp_exp_y2_21
      port map ( x => nY2,
                 r => nExpY2 );
  end generate;

  exp_y2_22 : if wF = 22 generate
    exp_y2 : fp_exp_exp_y2_22
      port map ( x => nY2,
                 r => nExpY2 );
  end generate;

  exp_y2_23 : if wF = 23 generate
    exp_y2 : fp_exp_exp_y2_23
      port map ( x => nY2,
                 r => nExpY2 );
  end generate;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library work;
use work.pkg_fp_exp.all;
use work.pkg_fp_exp_exp_y2.all;

entity fp_exp_exp_y2_clk is
  generic ( wF : positive );
  port ( nY2    : in  std_logic_vector(fp_exp_wy2(wF)-1 downto 0);
         nExpY2 : out std_logic_vector(fp_exp_wy2(wF) downto 0);
         clk    : in  std_logic );
end entity;

architecture arch of fp_exp_exp_y2_clk is
begin

  exp_y2_6 : if wF = 6 generate
    exp_y2 : fp_exp_exp_y2_6
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_7 : if wF = 7 generate
    exp_y2 : fp_exp_exp_y2_7
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_8 : if wF = 8 generate
    exp_y2 : fp_exp_exp_y2_8
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_9 : if wF = 9 generate
    exp_y2 : fp_exp_exp_y2_9
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_10 : if wF = 10 generate
    exp_y2 : fp_exp_exp_y2_10
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_11 : if wF = 11 generate
    exp_y2 : fp_exp_exp_y2_11
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_12 : if wF = 12 generate
    exp_y2 : fp_exp_exp_y2_12
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_13 : if wF = 13 generate
    exp_y2 : fp_exp_exp_y2_13
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_14 : if wF = 14 generate
    exp_y2 : fp_exp_exp_y2_14
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_15 : if wF = 15 generate
    exp_y2 : fp_exp_exp_y2_15
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_16 : if wF = 16 generate
    exp_y2 : fp_exp_exp_y2_16
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_17 : if wF = 17 generate
    exp_y2 : fp_exp_exp_y2_17
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_18 : if wF = 18 generate
    exp_y2 : fp_exp_exp_y2_18
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_19 : if wF = 19 generate
    exp_y2 : fp_exp_exp_y2_19
      port map ( nY2    => nY2,
                 nExpY2 => nExpY2(fp_exp_wy2(wF) downto 1) );
    nExpY2(0) <= '0';
  end generate;

  exp_y2_20 : if wF = 20 generate
    exp_y2 : fp_exp_exp_y2_20_clk
      port map ( x   => nY2,
                 r   => nExpY2,
                 clk => clk );
  end generate;

  exp_y2_21 : if wF = 21 generate
    exp_y2 : fp_exp_exp_y2_21_clk
      port map ( x   => nY2,
                 r   => nExpY2,
                 clk => clk );
  end generate;

  exp_y2_22 : if wF = 22 generate
    exp_y2 : fp_exp_exp_y2_22_clk
      port map ( x   => nY2,
                 r   => nExpY2,
                 clk => clk );
  end generate;

  exp_y2_23 : if wF = 23 generate
    exp_y2 : fp_exp_exp_y2_23_clk
      port map ( x   => nY2,
                 r   => nExpY2,
                 clk => clk );
  end generate;

end architecture;
