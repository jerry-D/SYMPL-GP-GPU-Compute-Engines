-- Copyright 2003-2006 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package pkg_fp_log_log is
  
  component fp_log_log_7 is
    port ( nX    : in  std_logic_vector(6 downto 0);
           nLogX : out std_logic_vector(8 downto 0) );
  end component;

  component fp_log_log_8 is
    port ( nX    : in  std_logic_vector(7 downto 0);
           nLogX : out std_logic_vector(9 downto 0) );
  end component;

  component fp_log_log_9 is
    port ( x : in  std_logic_vector(8 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component fp_log_log_10 is
    port ( x : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  component fp_log_log_11 is
    port ( x : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  component fp_log_log_11_clk is
    port ( x   : in  std_logic_vector(10 downto 0);
           r   : out std_logic_vector(13 downto 0);
           clk : in  std_logic );
  end component;

  component fp_log_log_12 is
    port ( x : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(15 downto 0) );
  end component;

  component fp_log_log_13 is
    port ( x : in  std_logic_vector(12 downto 0);
           r : out std_logic_vector(16 downto 0) );
  end component;

  component fp_log_log_14 is
    port ( x : in  std_logic_vector(13 downto 0);
           r : out std_logic_vector(16 downto 0) );
  end component;

  component fp_log_log_15 is
    port ( x : in  std_logic_vector(14 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

  component fp_log_log_16 is
    port ( x : in  std_logic_vector(15 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

  component fp_log_log_17 is
    port ( x : in  std_logic_vector(16 downto 0);
           r : out std_logic_vector(20 downto 0) );
  end component;

  component fp_log_log_18 is
    port ( x : in  std_logic_vector(17 downto 0);
           r : out std_logic_vector(21 downto 0) );
  end component;

  component fp_log_log_18_clk is
    port ( x   : in  std_logic_vector(17 downto 0);
           r   : out std_logic_vector(21 downto 0);
           clk : in  std_logic );
  end component;

  component fp_log_log_19 is
    port ( x : in  std_logic_vector(18 downto 0);
           r : out std_logic_vector(22 downto 0) );
  end component;

  component fp_log_log_20 is
    port ( x : in  std_logic_vector(19 downto 0);
           r : out std_logic_vector(23 downto 0) );
  end component;
  
  component fp_log_log_21 is
    port ( x : in  std_logic_vector(20 downto 0);
           r : out std_logic_vector(24 downto 0) );
  end component;

  component fp_log_log_22 is
    port ( x : in  std_logic_vector(21 downto 0);
           r : out std_logic_vector(25 downto 0) );
  end component;

  component fp_log_log_23 is
    port ( x : in  std_logic_vector(22 downto 0);
           r : out std_logic_vector(27 downto 0) );
  end component;

  component fp_log_log_24 is
    port ( x : in  std_logic_vector(23 downto 0);
           r : out std_logic_vector(28 downto 0) );
  end component;

  component fp_log_log_24_clk is
    port ( x   : in  std_logic_vector(23 downto 0);
           r   : out std_logic_vector(28 downto 0);
           clk : in  std_logic );
  end component;

end package;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_7 is
  port ( nX    : in  std_logic_vector(6 downto 0);
         nLogX : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of fp_log_log_7 is
begin

  with nX select
    nLogX <= "101100011" when "0000000", -- t[0] = 355
             "101100000" when "0000001", -- t[1] = 352
             "101011110" when "0000010", -- t[2] = 350
             "101011100" when "0000011", -- t[3] = 348
             "101011001" when "0000100", -- t[4] = 345
             "101010111" when "0000101", -- t[5] = 343
             "101010101" when "0000110", -- t[6] = 341
             "101010011" when "0000111", -- t[7] = 339
             "101010001" when "0001000", -- t[8] = 337
             "101001111" when "0001001", -- t[9] = 335
             "101001101" when "0001010", -- t[10] = 333
             "101001010" when "0001011", -- t[11] = 330
             "101001000" when "0001100", -- t[12] = 328
             "101000111" when "0001101", -- t[13] = 327
             "101000101" when "0001110", -- t[14] = 325
             "101000011" when "0001111", -- t[15] = 323
             "101000001" when "0010000", -- t[16] = 321
             "100111111" when "0010001", -- t[17] = 319
             "100111101" when "0010010", -- t[18] = 317
             "100111011" when "0010011", -- t[19] = 315
             "100111010" when "0010100", -- t[20] = 314
             "100111000" when "0010101", -- t[21] = 312
             "100110110" when "0010110", -- t[22] = 310
             "100110101" when "0010111", -- t[23] = 309
             "100110011" when "0011000", -- t[24] = 307
             "100110001" when "0011001", -- t[25] = 305
             "100110000" when "0011010", -- t[26] = 304
             "100101110" when "0011011", -- t[27] = 302
             "100101101" when "0011100", -- t[28] = 301
             "100101011" when "0011101", -- t[29] = 299
             "100101010" when "0011110", -- t[30] = 298
             "100101000" when "0011111", -- t[31] = 296
             "100100111" when "0100000", -- t[32] = 295
             "100100101" when "0100001", -- t[33] = 293
             "100100100" when "0100010", -- t[34] = 292
             "100100010" when "0100011", -- t[35] = 290
             "100100001" when "0100100", -- t[36] = 289
             "100100000" when "0100101", -- t[37] = 288
             "100011110" when "0100110", -- t[38] = 286
             "100011101" when "0100111", -- t[39] = 285
             "100011011" when "0101000", -- t[40] = 283
             "100011010" when "0101001", -- t[41] = 282
             "100011001" when "0101010", -- t[42] = 281
             "100011000" when "0101011", -- t[43] = 280
             "100010110" when "0101100", -- t[44] = 278
             "100010101" when "0101101", -- t[45] = 277
             "100010100" when "0101110", -- t[46] = 276
             "100010011" when "0101111", -- t[47] = 275
             "100010001" when "0110000", -- t[48] = 273
             "100010000" when "0110001", -- t[49] = 272
             "100001111" when "0110010", -- t[50] = 271
             "100001110" when "0110011", -- t[51] = 270
             "100001101" when "0110100", -- t[52] = 269
             "100001100" when "0110101", -- t[53] = 268
             "100001011" when "0110110", -- t[54] = 267
             "100001001" when "0110111", -- t[55] = 265
             "100001000" when "0111000", -- t[56] = 264
             "100000111" when "0111001", -- t[57] = 263
             "100000110" when "0111010", -- t[58] = 262
             "100000101" when "0111011", -- t[59] = 261
             "100000100" when "0111100", -- t[60] = 260
             "100000011" when "0111101", -- t[61] = 259
             "100000010" when "0111110", -- t[62] = 258
             "100000001" when "0111111", -- t[63] = 257
             "100000000" when "1000000", -- t[64] = 256
             "011111111" when "1000001", -- t[65] = 255
             "011111110" when "1000010", -- t[66] = 254
             "011111101" when "1000011", -- t[67] = 253
             "011111100" when "1000100", -- t[68] = 252
             "011111011" when "1000101", -- t[69] = 251
             "011111010" when "1000110", -- t[70] = 250
             "011111001" when "1000111", -- t[71] = 249
             "011111000" when "1001000", -- t[72] = 248
             "011110111" when "1001001", -- t[73] = 247
             "011110110" when "1001010", -- t[74] = 246
             "011110110" when "1001011", -- t[75] = 246
             "011110101" when "1001100", -- t[76] = 245
             "011110100" when "1001101", -- t[77] = 244
             "011110011" when "1001110", -- t[78] = 243
             "011110010" when "1001111", -- t[79] = 242
             "011110001" when "1010000", -- t[80] = 241
             "011110000" when "1010001", -- t[81] = 240
             "011110000" when "1010010", -- t[82] = 240
             "011101111" when "1010011", -- t[83] = 239
             "011101110" when "1010100", -- t[84] = 238
             "011101101" when "1010101", -- t[85] = 237
             "011101100" when "1010110", -- t[86] = 236
             "011101011" when "1010111", -- t[87] = 235
             "011101011" when "1011000", -- t[88] = 235
             "011101010" when "1011001", -- t[89] = 234
             "011101001" when "1011010", -- t[90] = 233
             "011101000" when "1011011", -- t[91] = 232
             "011101000" when "1011100", -- t[92] = 232
             "011100111" when "1011101", -- t[93] = 231
             "011100110" when "1011110", -- t[94] = 230
             "011100101" when "1011111", -- t[95] = 229
             "011100100" when "1100000", -- t[96] = 228
             "011100100" when "1100001", -- t[97] = 228
             "011100011" when "1100010", -- t[98] = 227
             "011100010" when "1100011", -- t[99] = 226
             "011100010" when "1100100", -- t[100] = 226
             "011100001" when "1100101", -- t[101] = 225
             "011100000" when "1100110", -- t[102] = 224
             "011011111" when "1100111", -- t[103] = 223
             "011011111" when "1101000", -- t[104] = 223
             "011011110" when "1101001", -- t[105] = 222
             "011011101" when "1101010", -- t[106] = 221
             "011011101" when "1101011", -- t[107] = 221
             "011011100" when "1101100", -- t[108] = 220
             "011011011" when "1101101", -- t[109] = 219
             "011011011" when "1101110", -- t[110] = 219
             "011011010" when "1101111", -- t[111] = 218
             "011011001" when "1110000", -- t[112] = 217
             "011011001" when "1110001", -- t[113] = 217
             "011011000" when "1110010", -- t[114] = 216
             "011010111" when "1110011", -- t[115] = 215
             "011010111" when "1110100", -- t[116] = 215
             "011010110" when "1110101", -- t[117] = 214
             "011010110" when "1110110", -- t[118] = 214
             "011010101" when "1110111", -- t[119] = 213
             "011010100" when "1111000", -- t[120] = 212
             "011010100" when "1111001", -- t[121] = 212
             "011010011" when "1111010", -- t[122] = 211
             "011010011" when "1111011", -- t[123] = 211
             "011010010" when "1111100", -- t[124] = 210
             "011010001" when "1111101", -- t[125] = 209
             "011010001" when "1111110", -- t[126] = 209
             "011010000" when "1111111", -- t[127] = 208
             "---------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_8 is
  port ( nX    : in  std_logic_vector(7 downto 0);
         nLogX : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of fp_log_log_8 is
begin

  with nX select
    nLogX <= "1011000110" when "00000000", -- t[0] = 710
             "1011000011" when "00000001", -- t[1] = 707
             "1011000001" when "00000010", -- t[2] = 705
             "1010111111" when "00000011", -- t[3] = 703
             "1010111100" when "00000100", -- t[4] = 700
             "1010111010" when "00000101", -- t[5] = 698
             "1010110111" when "00000110", -- t[6] = 695
             "1010110101" when "00000111", -- t[7] = 693
             "1010110011" when "00001000", -- t[8] = 691
             "1010110001" when "00001001", -- t[9] = 689
             "1010101110" when "00001010", -- t[10] = 686
             "1010101100" when "00001011", -- t[11] = 684
             "1010101010" when "00001100", -- t[12] = 682
             "1010101000" when "00001101", -- t[13] = 680
             "1010100110" when "00001110", -- t[14] = 678
             "1010100011" when "00001111", -- t[15] = 675
             "1010100001" when "00010000", -- t[16] = 673
             "1010011111" when "00010001", -- t[17] = 671
             "1010011101" when "00010010", -- t[18] = 669
             "1010011011" when "00010011", -- t[19] = 667
             "1010011001" when "00010100", -- t[20] = 665
             "1010010111" when "00010101", -- t[21] = 663
             "1010010101" when "00010110", -- t[22] = 661
             "1010010011" when "00010111", -- t[23] = 659
             "1010010001" when "00011000", -- t[24] = 657
             "1010001111" when "00011001", -- t[25] = 655
             "1010001101" when "00011010", -- t[26] = 653
             "1010001011" when "00011011", -- t[27] = 651
             "1010001001" when "00011100", -- t[28] = 649
             "1010000111" when "00011101", -- t[29] = 647
             "1010000101" when "00011110", -- t[30] = 645
             "1010000100" when "00011111", -- t[31] = 644
             "1010000010" when "00100000", -- t[32] = 642
             "1010000000" when "00100001", -- t[33] = 640
             "1001111110" when "00100010", -- t[34] = 638
             "1001111100" when "00100011", -- t[35] = 636
             "1001111010" when "00100100", -- t[36] = 634
             "1001111001" when "00100101", -- t[37] = 633
             "1001110111" when "00100110", -- t[38] = 631
             "1001110101" when "00100111", -- t[39] = 629
             "1001110011" when "00101000", -- t[40] = 627
             "1001110010" when "00101001", -- t[41] = 626
             "1001110000" when "00101010", -- t[42] = 624
             "1001101110" when "00101011", -- t[43] = 622
             "1001101101" when "00101100", -- t[44] = 621
             "1001101011" when "00101101", -- t[45] = 619
             "1001101001" when "00101110", -- t[46] = 617
             "1001101000" when "00101111", -- t[47] = 616
             "1001100110" when "00110000", -- t[48] = 614
             "1001100100" when "00110001", -- t[49] = 612
             "1001100011" when "00110010", -- t[50] = 611
             "1001100001" when "00110011", -- t[51] = 609
             "1001011111" when "00110100", -- t[52] = 607
             "1001011110" when "00110101", -- t[53] = 606
             "1001011100" when "00110110", -- t[54] = 604
             "1001011011" when "00110111", -- t[55] = 603
             "1001011001" when "00111000", -- t[56] = 601
             "1001011000" when "00111001", -- t[57] = 600
             "1001010110" when "00111010", -- t[58] = 598
             "1001010101" when "00111011", -- t[59] = 597
             "1001010011" when "00111100", -- t[60] = 595
             "1001010010" when "00111101", -- t[61] = 594
             "1001010000" when "00111110", -- t[62] = 592
             "1001001111" when "00111111", -- t[63] = 591
             "1001001101" when "01000000", -- t[64] = 589
             "1001001100" when "01000001", -- t[65] = 588
             "1001001010" when "01000010", -- t[66] = 586
             "1001001001" when "01000011", -- t[67] = 585
             "1001000111" when "01000100", -- t[68] = 583
             "1001000110" when "01000101", -- t[69] = 582
             "1001000101" when "01000110", -- t[70] = 581
             "1001000011" when "01000111", -- t[71] = 579
             "1001000010" when "01001000", -- t[72] = 578
             "1001000000" when "01001001", -- t[73] = 576
             "1000111111" when "01001010", -- t[74] = 575
             "1000111110" when "01001011", -- t[75] = 574
             "1000111100" when "01001100", -- t[76] = 572
             "1000111011" when "01001101", -- t[77] = 571
             "1000111010" when "01001110", -- t[78] = 570
             "1000111000" when "01001111", -- t[79] = 568
             "1000110111" when "01010000", -- t[80] = 567
             "1000110110" when "01010001", -- t[81] = 566
             "1000110100" when "01010010", -- t[82] = 564
             "1000110011" when "01010011", -- t[83] = 563
             "1000110010" when "01010100", -- t[84] = 562
             "1000110001" when "01010101", -- t[85] = 561
             "1000101111" when "01010110", -- t[86] = 559
             "1000101110" when "01010111", -- t[87] = 558
             "1000101101" when "01011000", -- t[88] = 557
             "1000101011" when "01011001", -- t[89] = 555
             "1000101010" when "01011010", -- t[90] = 554
             "1000101001" when "01011011", -- t[91] = 553
             "1000101000" when "01011100", -- t[92] = 552
             "1000100111" when "01011101", -- t[93] = 551
             "1000100101" when "01011110", -- t[94] = 549
             "1000100100" when "01011111", -- t[95] = 548
             "1000100011" when "01100000", -- t[96] = 547
             "1000100010" when "01100001", -- t[97] = 546
             "1000100001" when "01100010", -- t[98] = 545
             "1000011111" when "01100011", -- t[99] = 543
             "1000011110" when "01100100", -- t[100] = 542
             "1000011101" when "01100101", -- t[101] = 541
             "1000011100" when "01100110", -- t[102] = 540
             "1000011011" when "01100111", -- t[103] = 539
             "1000011010" when "01101000", -- t[104] = 538
             "1000011000" when "01101001", -- t[105] = 536
             "1000010111" when "01101010", -- t[106] = 535
             "1000010110" when "01101011", -- t[107] = 534
             "1000010101" when "01101100", -- t[108] = 533
             "1000010100" when "01101101", -- t[109] = 532
             "1000010011" when "01101110", -- t[110] = 531
             "1000010010" when "01101111", -- t[111] = 530
             "1000010001" when "01110000", -- t[112] = 529
             "1000010000" when "01110001", -- t[113] = 528
             "1000001111" when "01110010", -- t[114] = 527
             "1000001101" when "01110011", -- t[115] = 525
             "1000001100" when "01110100", -- t[116] = 524
             "1000001011" when "01110101", -- t[117] = 523
             "1000001010" when "01110110", -- t[118] = 522
             "1000001001" when "01110111", -- t[119] = 521
             "1000001000" when "01111000", -- t[120] = 520
             "1000000111" when "01111001", -- t[121] = 519
             "1000000110" when "01111010", -- t[122] = 518
             "1000000101" when "01111011", -- t[123] = 517
             "1000000100" when "01111100", -- t[124] = 516
             "1000000011" when "01111101", -- t[125] = 515
             "1000000010" when "01111110", -- t[126] = 514
             "1000000001" when "01111111", -- t[127] = 513
             "1000000000" when "10000000", -- t[128] = 512
             "0111111111" when "10000001", -- t[129] = 511
             "0111111110" when "10000010", -- t[130] = 510
             "0111111101" when "10000011", -- t[131] = 509
             "0111111100" when "10000100", -- t[132] = 508
             "0111111011" when "10000101", -- t[133] = 507
             "0111111010" when "10000110", -- t[134] = 506
             "0111111001" when "10000111", -- t[135] = 505
             "0111111000" when "10001000", -- t[136] = 504
             "0111110111" when "10001001", -- t[137] = 503
             "0111110110" when "10001010", -- t[138] = 502
             "0111110101" when "10001011", -- t[139] = 501
             "0111110100" when "10001100", -- t[140] = 500
             "0111110011" when "10001101", -- t[141] = 499
             "0111110010" when "10001110", -- t[142] = 498
             "0111110010" when "10001111", -- t[143] = 498
             "0111110001" when "10010000", -- t[144] = 497
             "0111110000" when "10010001", -- t[145] = 496
             "0111101111" when "10010010", -- t[146] = 495
             "0111101110" when "10010011", -- t[147] = 494
             "0111101101" when "10010100", -- t[148] = 493
             "0111101100" when "10010101", -- t[149] = 492
             "0111101011" when "10010110", -- t[150] = 491
             "0111101010" when "10010111", -- t[151] = 490
             "0111101001" when "10011000", -- t[152] = 489
             "0111101001" when "10011001", -- t[153] = 489
             "0111101000" when "10011010", -- t[154] = 488
             "0111100111" when "10011011", -- t[155] = 487
             "0111100110" when "10011100", -- t[156] = 486
             "0111100101" when "10011101", -- t[157] = 485
             "0111100100" when "10011110", -- t[158] = 484
             "0111100011" when "10011111", -- t[159] = 483
             "0111100010" when "10100000", -- t[160] = 482
             "0111100010" when "10100001", -- t[161] = 482
             "0111100001" when "10100010", -- t[162] = 481
             "0111100000" when "10100011", -- t[163] = 480
             "0111011111" when "10100100", -- t[164] = 479
             "0111011110" when "10100101", -- t[165] = 478
             "0111011101" when "10100110", -- t[166] = 477
             "0111011101" when "10100111", -- t[167] = 477
             "0111011100" when "10101000", -- t[168] = 476
             "0111011011" when "10101001", -- t[169] = 475
             "0111011010" when "10101010", -- t[170] = 474
             "0111011001" when "10101011", -- t[171] = 473
             "0111011000" when "10101100", -- t[172] = 472
             "0111011000" when "10101101", -- t[173] = 472
             "0111010111" when "10101110", -- t[174] = 471
             "0111010110" when "10101111", -- t[175] = 470
             "0111010101" when "10110000", -- t[176] = 469
             "0111010100" when "10110001", -- t[177] = 468
             "0111010100" when "10110010", -- t[178] = 468
             "0111010011" when "10110011", -- t[179] = 467
             "0111010010" when "10110100", -- t[180] = 466
             "0111010001" when "10110101", -- t[181] = 465
             "0111010001" when "10110110", -- t[182] = 465
             "0111010000" when "10110111", -- t[183] = 464
             "0111001111" when "10111000", -- t[184] = 463
             "0111001110" when "10111001", -- t[185] = 462
             "0111001101" when "10111010", -- t[186] = 461
             "0111001101" when "10111011", -- t[187] = 461
             "0111001100" when "10111100", -- t[188] = 460
             "0111001011" when "10111101", -- t[189] = 459
             "0111001010" when "10111110", -- t[190] = 458
             "0111001010" when "10111111", -- t[191] = 458
             "0111001001" when "11000000", -- t[192] = 457
             "0111001000" when "11000001", -- t[193] = 456
             "0111001000" when "11000010", -- t[194] = 456
             "0111000111" when "11000011", -- t[195] = 455
             "0111000110" when "11000100", -- t[196] = 454
             "0111000101" when "11000101", -- t[197] = 453
             "0111000101" when "11000110", -- t[198] = 453
             "0111000100" when "11000111", -- t[199] = 452
             "0111000011" when "11001000", -- t[200] = 451
             "0111000010" when "11001001", -- t[201] = 450
             "0111000010" when "11001010", -- t[202] = 450
             "0111000001" when "11001011", -- t[203] = 449
             "0111000000" when "11001100", -- t[204] = 448
             "0111000000" when "11001101", -- t[205] = 448
             "0110111111" when "11001110", -- t[206] = 447
             "0110111110" when "11001111", -- t[207] = 446
             "0110111110" when "11010000", -- t[208] = 446
             "0110111101" when "11010001", -- t[209] = 445
             "0110111100" when "11010010", -- t[210] = 444
             "0110111011" when "11010011", -- t[211] = 443
             "0110111011" when "11010100", -- t[212] = 443
             "0110111010" when "11010101", -- t[213] = 442
             "0110111001" when "11010110", -- t[214] = 441
             "0110111001" when "11010111", -- t[215] = 441
             "0110111000" when "11011000", -- t[216] = 440
             "0110110111" when "11011001", -- t[217] = 439
             "0110110111" when "11011010", -- t[218] = 439
             "0110110110" when "11011011", -- t[219] = 438
             "0110110101" when "11011100", -- t[220] = 437
             "0110110101" when "11011101", -- t[221] = 437
             "0110110100" when "11011110", -- t[222] = 436
             "0110110011" when "11011111", -- t[223] = 435
             "0110110011" when "11100000", -- t[224] = 435
             "0110110010" when "11100001", -- t[225] = 434
             "0110110001" when "11100010", -- t[226] = 433
             "0110110001" when "11100011", -- t[227] = 433
             "0110110000" when "11100100", -- t[228] = 432
             "0110110000" when "11100101", -- t[229] = 432
             "0110101111" when "11100110", -- t[230] = 431
             "0110101110" when "11100111", -- t[231] = 430
             "0110101110" when "11101000", -- t[232] = 430
             "0110101101" when "11101001", -- t[233] = 429
             "0110101100" when "11101010", -- t[234] = 428
             "0110101100" when "11101011", -- t[235] = 428
             "0110101011" when "11101100", -- t[236] = 427
             "0110101011" when "11101101", -- t[237] = 427
             "0110101010" when "11101110", -- t[238] = 426
             "0110101001" when "11101111", -- t[239] = 425
             "0110101001" when "11110000", -- t[240] = 425
             "0110101000" when "11110001", -- t[241] = 424
             "0110100111" when "11110010", -- t[242] = 423
             "0110100111" when "11110011", -- t[243] = 423
             "0110100110" when "11110100", -- t[244] = 422
             "0110100110" when "11110101", -- t[245] = 422
             "0110100101" when "11110110", -- t[246] = 421
             "0110100100" when "11110111", -- t[247] = 420
             "0110100100" when "11111000", -- t[248] = 420
             "0110100011" when "11111001", -- t[249] = 419
             "0110100011" when "11111010", -- t[250] = 419
             "0110100010" when "11111011", -- t[251] = 418
             "0110100010" when "11111100", -- t[252] = 418
             "0110100001" when "11111101", -- t[253] = 417
             "0110100000" when "11111110", -- t[254] = 416
             "0110100000" when "11111111", -- t[255] = 416
             "----------" when others;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 9; wO = 9.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 6; beta = 3;
--   T_0 (ROM):     alpha_0 = 6; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 4; beta_1 = 3.
-- Guard bits: g = 2.
-- Command line: logfp 9 9 1   rom 6 0   pm 4 3  ah 3 3 3  0 1  4 3 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 6; beta_0 = 0; wO_0 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_9_t0 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_9_t0 is
  signal x0   : std_logic_vector(5 downto 0);
  signal r0   : std_logic_vector(11 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "101100000111" when "000000", -- t[0] = 2823
          "101011100001" when "000001", -- t[1] = 2785
          "101010111100" when "000010", -- t[2] = 2748
          "101010011001" when "000011", -- t[3] = 2713
          "101001110111" when "000100", -- t[4] = 2679
          "101001010110" when "000101", -- t[5] = 2646
          "101000110111" when "000110", -- t[6] = 2615
          "101000011000" when "000111", -- t[7] = 2584
          "100111111011" when "001000", -- t[8] = 2555
          "100111011110" when "001001", -- t[9] = 2526
          "100111000010" when "001010", -- t[10] = 2498
          "100110100111" when "001011", -- t[11] = 2471
          "100110001101" when "001100", -- t[12] = 2445
          "100101110011" when "001101", -- t[13] = 2419
          "100101011011" when "001110", -- t[14] = 2395
          "100101000010" when "001111", -- t[15] = 2370
          "100100101011" when "010000", -- t[16] = 2347
          "100100010100" when "010001", -- t[17] = 2324
          "100011111110" when "010010", -- t[18] = 2302
          "100011101000" when "010011", -- t[19] = 2280
          "100011010011" when "010100", -- t[20] = 2259
          "100010111111" when "010101", -- t[21] = 2239
          "100010101011" when "010110", -- t[22] = 2219
          "100010010111" when "010111", -- t[23] = 2199
          "100010000100" when "011000", -- t[24] = 2180
          "100001110001" when "011001", -- t[25] = 2161
          "100001011111" when "011010", -- t[26] = 2143
          "100001001101" when "011011", -- t[27] = 2125
          "100000111100" when "011100", -- t[28] = 2108
          "100000101011" when "011101", -- t[29] = 2091
          "100000011010" when "011110", -- t[30] = 2074
          "100000001010" when "011111", -- t[31] = 2058
          "011111111010" when "100000", -- t[32] = 2042
          "011111101010" when "100001", -- t[33] = 2026
          "011111011010" when "100010", -- t[34] = 2010
          "011111001011" when "100011", -- t[35] = 1995
          "011110111101" when "100100", -- t[36] = 1981
          "011110101110" when "100101", -- t[37] = 1966
          "011110100000" when "100110", -- t[38] = 1952
          "011110010010" when "100111", -- t[39] = 1938
          "011110000100" when "101000", -- t[40] = 1924
          "011101110111" when "101001", -- t[41] = 1911
          "011101101010" when "101010", -- t[42] = 1898
          "011101011101" when "101011", -- t[43] = 1885
          "011101010000" when "101100", -- t[44] = 1872
          "011101000100" when "101101", -- t[45] = 1860
          "011100110111" when "101110", -- t[46] = 1847
          "011100101011" when "101111", -- t[47] = 1835
          "011100011111" when "110000", -- t[48] = 1823
          "011100010100" when "110001", -- t[49] = 1812
          "011100001000" when "110010", -- t[50] = 1800
          "011011111101" when "110011", -- t[51] = 1789
          "011011110010" when "110100", -- t[52] = 1778
          "011011100111" when "110101", -- t[53] = 1767
          "011011011100" when "110110", -- t[54] = 1756
          "011011010010" when "110111", -- t[55] = 1746
          "011011000111" when "111000", -- t[56] = 1735
          "011010111101" when "111001", -- t[57] = 1725
          "011010110011" when "111010", -- t[58] = 1715
          "011010101001" when "111011", -- t[59] = 1705
          "011010011111" when "111100", -- t[60] = 1695
          "011010010101" when "111101", -- t[61] = 1685
          "011010001100" when "111110", -- t[62] = 1676
          "011010000011" when "111111", -- t[63] = 1667
          "------------" when others;

  r(11 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 3; mu_1 = 3; lambda_1 = 3.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_9_t1_pow is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of fp_log_log_9_t1_pow is
  signal pp0 : std_logic_vector(1 downto 0);
  signal r0 : std_logic_vector(1 downto 0);
begin
  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(1 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 4; sigma'_1,1 = 2; wO_1,1 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_9_t1_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         s : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_log_log_9_t1_t1 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0010" when "000000", -- t[0] = 2
         "0110" when "000001", -- t[1] = 6
         "1011" when "000010", -- t[2] = 11
         "1111" when "000011", -- t[3] = 15
         "0001" when "000100", -- t[4] = 1
         "0101" when "000101", -- t[5] = 5
         "1001" when "000110", -- t[6] = 9
         "1101" when "000111", -- t[7] = 13
         "0001" when "001000", -- t[8] = 1
         "0101" when "001001", -- t[9] = 5
         "1000" when "001010", -- t[10] = 8
         "1100" when "001011", -- t[11] = 12
         "0001" when "001100", -- t[12] = 1
         "0100" when "001101", -- t[13] = 4
         "0111" when "001110", -- t[14] = 7
         "1010" when "001111", -- t[15] = 10
         "0001" when "010000", -- t[16] = 1
         "0100" when "010001", -- t[17] = 4
         "0110" when "010010", -- t[18] = 6
         "1001" when "010011", -- t[19] = 9
         "0001" when "010100", -- t[20] = 1
         "0011" when "010101", -- t[21] = 3
         "0110" when "010110", -- t[22] = 6
         "1000" when "010111", -- t[23] = 8
         "0001" when "011000", -- t[24] = 1
         "0011" when "011001", -- t[25] = 3
         "0101" when "011010", -- t[26] = 5
         "0111" when "011011", -- t[27] = 7
         "0001" when "011100", -- t[28] = 1
         "0011" when "011101", -- t[29] = 3
         "0101" when "011110", -- t[30] = 5
         "0111" when "011111", -- t[31] = 7
         "0000" when "100000", -- t[32] = 0
         "0010" when "100001", -- t[33] = 2
         "0100" when "100010", -- t[34] = 4
         "0110" when "100011", -- t[35] = 6
         "0000" when "100100", -- t[36] = 0
         "0010" when "100101", -- t[37] = 2
         "0100" when "100110", -- t[38] = 4
         "0110" when "100111", -- t[39] = 6
         "0000" when "101000", -- t[40] = 0
         "0010" when "101001", -- t[41] = 2
         "0100" when "101010", -- t[42] = 4
         "0101" when "101011", -- t[43] = 5
         "0000" when "101100", -- t[44] = 0
         "0010" when "101101", -- t[45] = 2
         "0011" when "101110", -- t[46] = 3
         "0101" when "101111", -- t[47] = 5
         "0000" when "110000", -- t[48] = 0
         "0010" when "110001", -- t[49] = 2
         "0011" when "110010", -- t[50] = 3
         "0101" when "110011", -- t[51] = 5
         "0000" when "110100", -- t[52] = 0
         "0010" when "110101", -- t[53] = 2
         "0011" when "110110", -- t[54] = 3
         "0100" when "110111", -- t[55] = 4
         "0000" when "111000", -- t[56] = 0
         "0001" when "111001", -- t[57] = 1
         "0011" when "111010", -- t[58] = 3
         "0100" when "111011", -- t[59] = 4
         "0000" when "111100", -- t[60] = 0
         "0001" when "111101", -- t[61] = 1
         "0010" when "111110", -- t[62] = 2
         "0100" when "111111", -- t[63] = 4
         "----" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 4; beta_1 = 3; lambda_1 = 3;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (ROM):  alpha_1,1 = 4; rho_1,1 = 0; sigma_1,1 = 3; wO_1,1 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_9_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         b : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_9_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(1 downto 0);
  signal s      : std_logic_vector(2 downto 0);
  component fp_log_log_9_t1_pow is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(2 downto 0) );
  end component;

  signal a_1    : std_logic_vector(3 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(1 downto 0);
  signal r0_1   : std_logic_vector(3 downto 0);
  signal r_1    : std_logic_vector(11 downto 0);
  component fp_log_log_9_t1_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;
begin
  sign <= not b(2);
  b0 <= b(1 downto 0) xor (1 downto 0 => sign);

  pow : fp_log_log_9_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(3 downto 0);
  sign_1 <= not s(2);
  s_1 <= s(1 downto 0) xor (1 downto 0 => sign_1);
  t_1 : fp_log_log_9_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_1 );
  r_1(3 downto 0) <=
    r0_1 xor (3 downto 0 => (not (sign xor sign_1)));
  r_1(11 downto 4) <= (11 downto 4 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_9 is
  port ( x : in  std_logic_vector(8 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_9 is
  signal a_0 : std_logic_vector(5 downto 0);
  signal r_0 : std_logic_vector(11 downto 0);
  component fp_log_log_9_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  signal a_1 : std_logic_vector(3 downto 0);
  signal b_1 : std_logic_vector(2 downto 0);
  signal r_1 : std_logic_vector(11 downto 0);
  component fp_log_log_9_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           b : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

begin
  a_0 <= x(8 downto 3);
  t_0 : fp_log_log_9_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(8 downto 5);
  b_1 <= x(2 downto 0);
  t_1 : fp_log_log_9_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  r <= r_0 + r_1;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 10; wO = 10.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 3;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 4; beta_1 = 3.
-- Guard bits: g = 3.
-- Command line: logfp 10 10 1   rom 7 0   pm 4 3  ah 3 3 3  0 1  4 3 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 14.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_10_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_10_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(13 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110000111011" when "0000000", -- t[0] = 11323
          "10101111101110" when "0000001", -- t[1] = 11246
          "10101110100010" when "0000010", -- t[2] = 11170
          "10101101011000" when "0000011", -- t[3] = 11096
          "10101100001111" when "0000100", -- t[4] = 11023
          "10101011000111" when "0000101", -- t[5] = 10951
          "10101010000001" when "0000110", -- t[6] = 10881
          "10101000111100" when "0000111", -- t[7] = 10812
          "10100111111001" when "0001000", -- t[8] = 10745
          "10100110110110" when "0001001", -- t[9] = 10678
          "10100101110100" when "0001010", -- t[10] = 10612
          "10100100110100" when "0001011", -- t[11] = 10548
          "10100011110101" when "0001100", -- t[12] = 10485
          "10100010110111" when "0001101", -- t[13] = 10423
          "10100001111010" when "0001110", -- t[14] = 10362
          "10100000111101" when "0001111", -- t[15] = 10301
          "10100000000010" when "0010000", -- t[16] = 10242
          "10011111001000" when "0010001", -- t[17] = 10184
          "10011110001110" when "0010010", -- t[18] = 10126
          "10011101010110" when "0010011", -- t[19] = 10070
          "10011100011110" when "0010100", -- t[20] = 10014
          "10011011101000" when "0010101", -- t[21] = 9960
          "10011010110010" when "0010110", -- t[22] = 9906
          "10011001111100" when "0010111", -- t[23] = 9852
          "10011001001000" when "0011000", -- t[24] = 9800
          "10011000010100" when "0011001", -- t[25] = 9748
          "10010111100010" when "0011010", -- t[26] = 9698
          "10010110101111" when "0011011", -- t[27] = 9647
          "10010101111110" when "0011100", -- t[28] = 9598
          "10010101001101" when "0011101", -- t[29] = 9549
          "10010100011101" when "0011110", -- t[30] = 9501
          "10010011101110" when "0011111", -- t[31] = 9454
          "10010010111111" when "0100000", -- t[32] = 9407
          "10010010010001" when "0100001", -- t[33] = 9361
          "10010001100011" when "0100010", -- t[34] = 9315
          "10010000110110" when "0100011", -- t[35] = 9270
          "10010000001010" when "0100100", -- t[36] = 9226
          "10001111011110" when "0100101", -- t[37] = 9182
          "10001110110011" when "0100110", -- t[38] = 9139
          "10001110001000" when "0100111", -- t[39] = 9096
          "10001101011110" when "0101000", -- t[40] = 9054
          "10001100110100" when "0101001", -- t[41] = 9012
          "10001100001011" when "0101010", -- t[42] = 8971
          "10001011100011" when "0101011", -- t[43] = 8931
          "10001010111011" when "0101100", -- t[44] = 8891
          "10001010010011" when "0101101", -- t[45] = 8851
          "10001001101100" when "0101110", -- t[46] = 8812
          "10001001000101" when "0101111", -- t[47] = 8773
          "10001000011111" when "0110000", -- t[48] = 8735
          "10000111111001" when "0110001", -- t[49] = 8697
          "10000111010100" when "0110010", -- t[50] = 8660
          "10000110101111" when "0110011", -- t[51] = 8623
          "10000110001010" when "0110100", -- t[52] = 8586
          "10000101100110" when "0110101", -- t[53] = 8550
          "10000101000011" when "0110110", -- t[54] = 8515
          "10000100011111" when "0110111", -- t[55] = 8479
          "10000011111100" when "0111000", -- t[56] = 8444
          "10000011011010" when "0111001", -- t[57] = 8410
          "10000010111000" when "0111010", -- t[58] = 8376
          "10000010010110" when "0111011", -- t[59] = 8342
          "10000001110101" when "0111100", -- t[60] = 8309
          "10000001010100" when "0111101", -- t[61] = 8276
          "10000000110011" when "0111110", -- t[62] = 8243
          "10000000010011" when "0111111", -- t[63] = 8211
          "01111111110011" when "1000000", -- t[64] = 8179
          "01111111010011" when "1000001", -- t[65] = 8147
          "01111110110011" when "1000010", -- t[66] = 8115
          "01111110010100" when "1000011", -- t[67] = 8084
          "01111101110110" when "1000100", -- t[68] = 8054
          "01111101010111" when "1000101", -- t[69] = 8023
          "01111100111001" when "1000110", -- t[70] = 7993
          "01111100011011" when "1000111", -- t[71] = 7963
          "01111011111110" when "1001000", -- t[72] = 7934
          "01111011100001" when "1001001", -- t[73] = 7905
          "01111011000100" when "1001010", -- t[74] = 7876
          "01111010100111" when "1001011", -- t[75] = 7847
          "01111010001011" when "1001100", -- t[76] = 7819
          "01111001101110" when "1001101", -- t[77] = 7790
          "01111001010011" when "1001110", -- t[78] = 7763
          "01111000110111" when "1001111", -- t[79] = 7735
          "01111000011100" when "1010000", -- t[80] = 7708
          "01111000000001" when "1010001", -- t[81] = 7681
          "01110111100110" when "1010010", -- t[82] = 7654
          "01110111001011" when "1010011", -- t[83] = 7627
          "01110110110001" when "1010100", -- t[84] = 7601
          "01110110010111" when "1010101", -- t[85] = 7575
          "01110101111101" when "1010110", -- t[86] = 7549
          "01110101100011" when "1010111", -- t[87] = 7523
          "01110101001010" when "1011000", -- t[88] = 7498
          "01110100110000" when "1011001", -- t[89] = 7472
          "01110100011000" when "1011010", -- t[90] = 7448
          "01110011111111" when "1011011", -- t[91] = 7423
          "01110011100110" when "1011100", -- t[92] = 7398
          "01110011001110" when "1011101", -- t[93] = 7374
          "01110010110110" when "1011110", -- t[94] = 7350
          "01110010011110" when "1011111", -- t[95] = 7326
          "01110010000110" when "1100000", -- t[96] = 7302
          "01110001101111" when "1100001", -- t[97] = 7279
          "01110001010111" when "1100010", -- t[98] = 7255
          "01110001000000" when "1100011", -- t[99] = 7232
          "01110000101001" when "1100100", -- t[100] = 7209
          "01110000010011" when "1100101", -- t[101] = 7187
          "01101111111100" when "1100110", -- t[102] = 7164
          "01101111100110" when "1100111", -- t[103] = 7142
          "01101111001111" when "1101000", -- t[104] = 7119
          "01101110111001" when "1101001", -- t[105] = 7097
          "01101110100100" when "1101010", -- t[106] = 7076
          "01101110001110" when "1101011", -- t[107] = 7054
          "01101101111000" when "1101100", -- t[108] = 7032
          "01101101100011" when "1101101", -- t[109] = 7011
          "01101101001110" when "1101110", -- t[110] = 6990
          "01101100111001" when "1101111", -- t[111] = 6969
          "01101100100100" when "1110000", -- t[112] = 6948
          "01101100001111" when "1110001", -- t[113] = 6927
          "01101011111011" when "1110010", -- t[114] = 6907
          "01101011100111" when "1110011", -- t[115] = 6887
          "01101011010010" when "1110100", -- t[116] = 6866
          "01101010111110" when "1110101", -- t[117] = 6846
          "01101010101011" when "1110110", -- t[118] = 6827
          "01101010010111" when "1110111", -- t[119] = 6807
          "01101010000011" when "1111000", -- t[120] = 6787
          "01101001110000" when "1111001", -- t[121] = 6768
          "01101001011100" when "1111010", -- t[122] = 6748
          "01101001001001" when "1111011", -- t[123] = 6729
          "01101000110110" when "1111100", -- t[124] = 6710
          "01101000100011" when "1111101", -- t[125] = 6691
          "01101000010001" when "1111110", -- t[126] = 6673
          "01100111111110" when "1111111", -- t[127] = 6654
          "--------------" when others;

  r(13 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 3; mu_1 = 3; lambda_1 = 3.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_10_t1_pow is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of fp_log_log_10_t1_pow is
  signal pp0 : std_logic_vector(1 downto 0);
  signal r0 : std_logic_vector(1 downto 0);
begin
  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(1 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 4; sigma'_1,1 = 2; wO_1,1 = 5.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_10_t1_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         s : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of fp_log_log_10_t1_t1 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a & s;

  with x select
    r <= "00100" when "000000", -- t[0] = 4
         "01101" when "000001", -- t[1] = 13
         "10110" when "000010", -- t[2] = 22
         "11111" when "000011", -- t[3] = 31
         "00011" when "000100", -- t[4] = 3
         "01011" when "000101", -- t[5] = 11
         "10011" when "000110", -- t[6] = 19
         "11011" when "000111", -- t[7] = 27
         "00011" when "001000", -- t[8] = 3
         "01010" when "001001", -- t[9] = 10
         "10001" when "001010", -- t[10] = 17
         "11000" when "001011", -- t[11] = 24
         "00011" when "001100", -- t[12] = 3
         "01001" when "001101", -- t[13] = 9
         "01111" when "001110", -- t[14] = 15
         "10101" when "001111", -- t[15] = 21
         "00010" when "010000", -- t[16] = 2
         "01000" when "010001", -- t[17] = 8
         "01101" when "010010", -- t[18] = 13
         "10011" when "010011", -- t[19] = 19
         "00010" when "010100", -- t[20] = 2
         "00111" when "010101", -- t[21] = 7
         "01100" when "010110", -- t[22] = 12
         "10001" when "010111", -- t[23] = 17
         "00010" when "011000", -- t[24] = 2
         "00110" when "011001", -- t[25] = 6
         "01011" when "011010", -- t[26] = 11
         "01111" when "011011", -- t[27] = 15
         "00010" when "011100", -- t[28] = 2
         "00110" when "011101", -- t[29] = 6
         "01010" when "011110", -- t[30] = 10
         "01110" when "011111", -- t[31] = 14
         "00001" when "100000", -- t[32] = 1
         "00101" when "100001", -- t[33] = 5
         "01001" when "100010", -- t[34] = 9
         "01101" when "100011", -- t[35] = 13
         "00001" when "100100", -- t[36] = 1
         "00101" when "100101", -- t[37] = 5
         "01000" when "100110", -- t[38] = 8
         "01100" when "100111", -- t[39] = 12
         "00001" when "101000", -- t[40] = 1
         "00100" when "101001", -- t[41] = 4
         "01000" when "101010", -- t[42] = 8
         "01011" when "101011", -- t[43] = 11
         "00001" when "101100", -- t[44] = 1
         "00100" when "101101", -- t[45] = 4
         "00111" when "101110", -- t[46] = 7
         "01010" when "101111", -- t[47] = 10
         "00001" when "110000", -- t[48] = 1
         "00100" when "110001", -- t[49] = 4
         "00111" when "110010", -- t[50] = 7
         "01010" when "110011", -- t[51] = 10
         "00001" when "110100", -- t[52] = 1
         "00100" when "110101", -- t[53] = 4
         "00110" when "110110", -- t[54] = 6
         "01001" when "110111", -- t[55] = 9
         "00001" when "111000", -- t[56] = 1
         "00011" when "111001", -- t[57] = 3
         "00110" when "111010", -- t[58] = 6
         "01000" when "111011", -- t[59] = 8
         "00001" when "111100", -- t[60] = 1
         "00011" when "111101", -- t[61] = 3
         "00101" when "111110", -- t[62] = 5
         "01000" when "111111", -- t[63] = 8
         "-----" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 4; beta_1 = 3; lambda_1 = 3;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (ROM):  alpha_1,1 = 4; rho_1,1 = 0; sigma_1,1 = 3; wO_1,1 = 5.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_10_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         b : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_10_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(1 downto 0);
  signal s      : std_logic_vector(2 downto 0);
  component fp_log_log_10_t1_pow is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(2 downto 0) );
  end component;

  signal a_1    : std_logic_vector(3 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(1 downto 0);
  signal r0_1   : std_logic_vector(4 downto 0);
  signal r_1    : std_logic_vector(13 downto 0);
  component fp_log_log_10_t1_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;
begin
  sign <= not b(2);
  b0 <= b(1 downto 0) xor (1 downto 0 => sign);

  pow : fp_log_log_10_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(3 downto 0);
  sign_1 <= not s(2);
  s_1 <= s(1 downto 0) xor (1 downto 0 => sign_1);
  t_1 : fp_log_log_10_t1_t1
    port map ( a => a_1,
               s => s_1,
               r => r0_1 );
  r_1(4 downto 0) <=
    r0_1 xor (4 downto 0 => (not (sign xor sign_1)));
  r_1(13 downto 5) <= (13 downto 5 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_10 is
  port ( x : in  std_logic_vector(9 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_10 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(13 downto 0);
  component fp_log_log_10_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1 : std_logic_vector(3 downto 0);
  signal b_1 : std_logic_vector(2 downto 0);
  signal r_1 : std_logic_vector(13 downto 0);
  component fp_log_log_10_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           b : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

begin
  a_0 <= x(9 downto 3);
  t_0 : fp_log_log_10_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(9 downto 6);
  b_1 <= x(2 downto 0);
  t_1 : fp_log_log_10_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  r <= r_0 + r_1;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 11; wO = 11.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 4;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 5; beta_1 = 4.
-- Guard bits: g = 2.
-- Command line: logfp 11 11 1   rom 7 0   pm 5 4  ah 4 4 4  1 0  5 4 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 14.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_11_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_11_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(13 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110000111000" when "0000000", -- t[0] = 11320
          "10101111101011" when "0000001", -- t[1] = 11243
          "10101110100000" when "0000010", -- t[2] = 11168
          "10101101010110" when "0000011", -- t[3] = 11094
          "10101100001101" when "0000100", -- t[4] = 11021
          "10101011000101" when "0000101", -- t[5] = 10949
          "10101001111111" when "0000110", -- t[6] = 10879
          "10101000111010" when "0000111", -- t[7] = 10810
          "10100111110110" when "0001000", -- t[8] = 10742
          "10100110110100" when "0001001", -- t[9] = 10676
          "10100101110010" when "0001010", -- t[10] = 10610
          "10100100110010" when "0001011", -- t[11] = 10546
          "10100011110011" when "0001100", -- t[12] = 10483
          "10100010110101" when "0001101", -- t[13] = 10421
          "10100001111000" when "0001110", -- t[14] = 10360
          "10100000111100" when "0001111", -- t[15] = 10300
          "10100000000000" when "0010000", -- t[16] = 10240
          "10011111000110" when "0010001", -- t[17] = 10182
          "10011110001101" when "0010010", -- t[18] = 10125
          "10011101010100" when "0010011", -- t[19] = 10068
          "10011100011101" when "0010100", -- t[20] = 10013
          "10011011100110" when "0010101", -- t[21] = 9958
          "10011010110000" when "0010110", -- t[22] = 9904
          "10011001111011" when "0010111", -- t[23] = 9851
          "10011001000110" when "0011000", -- t[24] = 9798
          "10011000010011" when "0011001", -- t[25] = 9747
          "10010111100000" when "0011010", -- t[26] = 9696
          "10010110101110" when "0011011", -- t[27] = 9646
          "10010101111100" when "0011100", -- t[28] = 9596
          "10010101001100" when "0011101", -- t[29] = 9548
          "10010100011100" when "0011110", -- t[30] = 9500
          "10010011101100" when "0011111", -- t[31] = 9452
          "10010010111101" when "0100000", -- t[32] = 9405
          "10010010001111" when "0100001", -- t[33] = 9359
          "10010001100010" when "0100010", -- t[34] = 9314
          "10010000110101" when "0100011", -- t[35] = 9269
          "10010000001001" when "0100100", -- t[36] = 9225
          "10001111011101" when "0100101", -- t[37] = 9181
          "10001110110010" when "0100110", -- t[38] = 9138
          "10001110000111" when "0100111", -- t[39] = 9095
          "10001101011101" when "0101000", -- t[40] = 9053
          "10001100110011" when "0101001", -- t[41] = 9011
          "10001100001010" when "0101010", -- t[42] = 8970
          "10001011100001" when "0101011", -- t[43] = 8929
          "10001010111001" when "0101100", -- t[44] = 8889
          "10001010010010" when "0101101", -- t[45] = 8850
          "10001001101011" when "0101110", -- t[46] = 8811
          "10001001000100" when "0101111", -- t[47] = 8772
          "10001000011110" when "0110000", -- t[48] = 8734
          "10000111111000" when "0110001", -- t[49] = 8696
          "10000111010011" when "0110010", -- t[50] = 8659
          "10000110101110" when "0110011", -- t[51] = 8622
          "10000110001001" when "0110100", -- t[52] = 8585
          "10000101100101" when "0110101", -- t[53] = 8549
          "10000101000010" when "0110110", -- t[54] = 8514
          "10000100011110" when "0110111", -- t[55] = 8478
          "10000011111011" when "0111000", -- t[56] = 8443
          "10000011011001" when "0111001", -- t[57] = 8409
          "10000010110111" when "0111010", -- t[58] = 8375
          "10000010010101" when "0111011", -- t[59] = 8341
          "10000001110100" when "0111100", -- t[60] = 8308
          "10000001010011" when "0111101", -- t[61] = 8275
          "10000000110010" when "0111110", -- t[62] = 8242
          "10000000010010" when "0111111", -- t[63] = 8210
          "01111111110010" when "1000000", -- t[64] = 8178
          "01111111010010" when "1000001", -- t[65] = 8146
          "01111110110011" when "1000010", -- t[66] = 8115
          "01111110010011" when "1000011", -- t[67] = 8083
          "01111101110101" when "1000100", -- t[68] = 8053
          "01111101010110" when "1000101", -- t[69] = 8022
          "01111100111000" when "1000110", -- t[70] = 7992
          "01111100011010" when "1000111", -- t[71] = 7962
          "01111011111101" when "1001000", -- t[72] = 7933
          "01111011100000" when "1001001", -- t[73] = 7904
          "01111011000011" when "1001010", -- t[74] = 7875
          "01111010100110" when "1001011", -- t[75] = 7846
          "01111010001010" when "1001100", -- t[76] = 7818
          "01111001101110" when "1001101", -- t[77] = 7790
          "01111001010010" when "1001110", -- t[78] = 7762
          "01111000110110" when "1001111", -- t[79] = 7734
          "01111000011011" when "1010000", -- t[80] = 7707
          "01111000000000" when "1010001", -- t[81] = 7680
          "01110111100101" when "1010010", -- t[82] = 7653
          "01110111001010" when "1010011", -- t[83] = 7626
          "01110110110000" when "1010100", -- t[84] = 7600
          "01110110010110" when "1010101", -- t[85] = 7574
          "01110101111100" when "1010110", -- t[86] = 7548
          "01110101100010" when "1010111", -- t[87] = 7522
          "01110101001001" when "1011000", -- t[88] = 7497
          "01110100110000" when "1011001", -- t[89] = 7472
          "01110100010111" when "1011010", -- t[90] = 7447
          "01110011111110" when "1011011", -- t[91] = 7422
          "01110011100101" when "1011100", -- t[92] = 7397
          "01110011001101" when "1011101", -- t[93] = 7373
          "01110010110101" when "1011110", -- t[94] = 7349
          "01110010011101" when "1011111", -- t[95] = 7325
          "01110010000101" when "1100000", -- t[96] = 7301
          "01110001101110" when "1100001", -- t[97] = 7278
          "01110001010111" when "1100010", -- t[98] = 7255
          "01110000111111" when "1100011", -- t[99] = 7231
          "01110000101001" when "1100100", -- t[100] = 7209
          "01110000010010" when "1100101", -- t[101] = 7186
          "01101111111011" when "1100110", -- t[102] = 7163
          "01101111100101" when "1100111", -- t[103] = 7141
          "01101111001111" when "1101000", -- t[104] = 7119
          "01101110111001" when "1101001", -- t[105] = 7097
          "01101110100011" when "1101010", -- t[106] = 7075
          "01101110001101" when "1101011", -- t[107] = 7053
          "01101101111000" when "1101100", -- t[108] = 7032
          "01101101100010" when "1101101", -- t[109] = 7010
          "01101101001101" when "1101110", -- t[110] = 6989
          "01101100111000" when "1101111", -- t[111] = 6968
          "01101100100011" when "1110000", -- t[112] = 6947
          "01101100001111" when "1110001", -- t[113] = 6927
          "01101011111010" when "1110010", -- t[114] = 6906
          "01101011100110" when "1110011", -- t[115] = 6886
          "01101011010010" when "1110100", -- t[116] = 6866
          "01101010111110" when "1110101", -- t[117] = 6846
          "01101010101010" when "1110110", -- t[118] = 6826
          "01101010010110" when "1110111", -- t[119] = 6806
          "01101010000011" when "1111000", -- t[120] = 6787
          "01101001101111" when "1111001", -- t[121] = 6767
          "01101001011100" when "1111010", -- t[122] = 6748
          "01101001001001" when "1111011", -- t[123] = 6729
          "01101000110110" when "1111100", -- t[124] = 6710
          "01101000100011" when "1111101", -- t[125] = 6691
          "01101000010000" when "1111110", -- t[126] = 6672
          "01100111111101" when "1111111", -- t[127] = 6653
          "--------------" when others;

  r(13 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 4; mu_1 = 4; lambda_1 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_11_t1_pow is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_log_log_11_t1_pow is
  signal pp0 : std_logic_vector(2 downto 0);
  signal r0 : std_logic_vector(2 downto 0);
begin
  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(2 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 5; wO_1,1 = 7.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_11_t1_t1 is
  port ( a : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_log_log_11_t1_t1 is
  signal x : std_logic_vector(4 downto 0);
begin
  x <= a;

  with x select
    r <= "1001100" when "00000", -- t[0] = 76
         "1000110" when "00001", -- t[1] = 70
         "1000001" when "00010", -- t[2] = 65
         "0111101" when "00011", -- t[3] = 61
         "0111001" when "00100", -- t[4] = 57
         "0110110" when "00101", -- t[5] = 54
         "0110011" when "00110", -- t[6] = 51
         "0110000" when "00111", -- t[7] = 48
         "0101110" when "01000", -- t[8] = 46
         "0101011" when "01001", -- t[9] = 43
         "0101001" when "01010", -- t[10] = 41
         "0100111" when "01011", -- t[11] = 39
         "0100101" when "01100", -- t[12] = 37
         "0100100" when "01101", -- t[13] = 36
         "0100010" when "01110", -- t[14] = 34
         "0100001" when "01111", -- t[15] = 33
         "0011111" when "10000", -- t[16] = 31
         "0011110" when "10001", -- t[17] = 30
         "0011101" when "10010", -- t[18] = 29
         "0011100" when "10011", -- t[19] = 28
         "0011011" when "10100", -- t[20] = 27
         "0011010" when "10101", -- t[21] = 26
         "0011001" when "10110", -- t[22] = 25
         "0011000" when "10111", -- t[23] = 24
         "0010111" when "11000", -- t[24] = 23
         "0010111" when "11001", -- t[25] = 23
         "0010110" when "11010", -- t[26] = 22
         "0010101" when "11011", -- t[27] = 21
         "0010100" when "11100", -- t[28] = 20
         "0010100" when "11101", -- t[29] = 20
         "0010011" when "11110", -- t[30] = 19
         "0010011" when "11111", -- t[31] = 19
         "-------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 5; beta_1 = 4; lambda_1 = 4;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 5; rho_1,1 = 0; sigma_1,1 = 4; wO_1,1 = 7.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_11_t1 is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_11_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(2 downto 0);
  signal s      : std_logic_vector(3 downto 0);
  component fp_log_log_11_t1_pow is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  signal a_1    : std_logic_vector(4 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(2 downto 0);
  signal k_1    : std_logic_vector(6 downto 0);
  signal r0_1   : std_logic_vector(11 downto 0);
  signal r_1    : std_logic_vector(13 downto 0);
  component fp_log_log_11_t1_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;
begin
  sign <= not b(3);
  b0 <= b(2 downto 0) xor (2 downto 0 => sign);

  pow : fp_log_log_11_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(4 downto 0);
  sign_1 <= not s(3);
  s_1 <= s(2 downto 0) xor (2 downto 0 => sign_1);
  t_1 : fp_log_log_11_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(6 downto 0) <=
    r0_1(11 downto 5) xor (11 downto 5 => (not (sign xor sign_1)));
  r_1(13 downto 7) <= (13 downto 7 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_11_t1_clk is
  port ( a   : in  std_logic_vector(4 downto 0);
         b   : in  std_logic_vector(3 downto 0);
         r   : out std_logic_vector(13 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_11_t1_clk is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(2 downto 0);
  signal s      : std_logic_vector(3 downto 0);
  component fp_log_log_11_t1_pow is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  signal a_1     : std_logic_vector(4 downto 0);
  signal sign_1  : std_logic;
  signal sgn_1_0 : std_logic;
  signal sgn_1   : std_logic;
  signal s_1_0   : std_logic_vector(2 downto 0);
  signal s_1     : std_logic_vector(2 downto 0);
  signal k_1_0   : std_logic_vector(6 downto 0);
  signal k_1     : std_logic_vector(6 downto 0);
  signal r0_1    : std_logic_vector(11 downto 0);
  signal r_1     : std_logic_vector(13 downto 0);
  component fp_log_log_11_t1_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;
begin
  sign <= not b(3);
  b0 <= b(2 downto 0) xor (2 downto 0 => sign);

  pow : fp_log_log_11_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(4 downto 0);
  sign_1 <= not s(3);
  sgn_1_0 <= sign xor sign_1;
  s_1_0 <= s(2 downto 0) xor (2 downto 0 => sign_1);
  t_1 : fp_log_log_11_t1_t1
    port map ( a => a_1,
               r => k_1_0 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(6 downto 0) <=
    r0_1(11 downto 5) xor (11 downto 5 => (not (sgn_1)));
  r_1(13 downto 7) <= (13 downto 7 => (not (sgn_1)));

  process(clk)
  begin
    if clk'event and clk = '1' then
      sgn_1 <= sgn_1_0;
      s_1   <= s_1_0;
      k_1   <= k_1_0;
    end if;
  end process;

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_11 is
  port ( x : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_11 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(13 downto 0);
  component fp_log_log_11_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1 : std_logic_vector(4 downto 0);
  signal b_1 : std_logic_vector(3 downto 0);
  signal r_1 : std_logic_vector(13 downto 0);
  component fp_log_log_11_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

begin
  a_0 <= x(10 downto 4);
  t_0 : fp_log_log_11_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(10 downto 6);
  b_1 <= x(3 downto 0);
  t_1 : fp_log_log_11_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  r <= r_0 + r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_11_clk is
  port ( x   : in  std_logic_vector(10 downto 0);
         r   : out std_logic_vector(13 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_11_clk is
  signal a_0_0 : std_logic_vector(6 downto 0);
  signal a_0   : std_logic_vector(6 downto 0);
  signal r_0   : std_logic_vector(13 downto 0);
  component fp_log_log_11_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1   : std_logic_vector(4 downto 0);
  signal b_1   : std_logic_vector(3 downto 0);
  signal r_1   : std_logic_vector(13 downto 0);
  component fp_log_log_11_t1_clk is
    port ( a   : in  std_logic_vector(4 downto 0);
           b   : in  std_logic_vector(3 downto 0);
           r   : out std_logic_vector(13 downto 0);
           clk : in  std_logic );
  end component;

begin
  a_0_0 <= x(10 downto 4);
  t_0 : fp_log_log_11_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(10 downto 6);
  b_1 <= x(3 downto 0);
  t_1 : fp_log_log_11_t1_clk
    port map ( a   => a_1,
               b   => b_1,
               r   => r_1,
               clk => clk );

  process(clk)
  begin
    if clk'event and clk = '1' then
      a_0 <= a_0_0;
    end if;
  end process;

  r <= r_0 + r_1;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 12; wO = 12.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 6; beta = 6;
--   T_0 (ROM):     alpha_0 = 6; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 6; beta_1 = 6.
-- Guard bits: g = 3.
-- Command line: logfp 12 12 1   rom 6 0   pm 6 6  ah 6 6 6  1 1  6 4 0  4 2 4


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 6; beta_0 = 0; wO_0 = 16.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_12_t0 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of fp_log_log_12_t0 is
  signal x0   : std_logic_vector(5 downto 0);
  signal r0   : std_logic_vector(15 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "1011000001000010" when "000000", -- t[0] = 45122
          "1010110111100101" when "000001", -- t[1] = 44517
          "1010101110011111" when "000010", -- t[2] = 43935
          "1010100101101101" when "000011", -- t[3] = 43373
          "1010011101010000" when "000100", -- t[4] = 42832
          "1010010101000101" when "000101", -- t[5] = 42309
          "1010001101001011" when "000110", -- t[6] = 41803
          "1010000101100010" when "000111", -- t[7] = 41314
          "1001111110001000" when "001000", -- t[8] = 40840
          "1001110110111110" when "001001", -- t[9] = 40382
          "1001110000000001" when "001010", -- t[10] = 39937
          "1001101001010001" when "001011", -- t[11] = 39505
          "1001100010101111" when "001100", -- t[12] = 39087
          "1001011100011000" when "001101", -- t[13] = 38680
          "1001010110001100" when "001110", -- t[14] = 38284
          "1001010000001100" when "001111", -- t[15] = 37900
          "1001001010010110" when "010000", -- t[16] = 37526
          "1001000100101010" when "010001", -- t[17] = 37162
          "1000111111000111" when "010010", -- t[18] = 36807
          "1000111001101101" when "010011", -- t[19] = 36461
          "1000110100011100" when "010100", -- t[20] = 36124
          "1000101111010100" when "010101", -- t[21] = 35796
          "1000101010010011" when "010110", -- t[22] = 35475
          "1000100101011010" when "010111", -- t[23] = 35162
          "1000100000101000" when "011000", -- t[24] = 34856
          "1000011011111110" when "011001", -- t[25] = 34558
          "1000010111011010" when "011010", -- t[26] = 34266
          "1000010010111101" when "011011", -- t[27] = 33981
          "1000001110100110" when "011100", -- t[28] = 33702
          "1000001010010101" when "011101", -- t[29] = 33429
          "1000000110001010" when "011110", -- t[30] = 33162
          "1000000010000100" when "011111", -- t[31] = 32900
          "0111111110000100" when "100000", -- t[32] = 32644
          "0111111010001001" when "100001", -- t[33] = 32393
          "0111110110010011" when "100010", -- t[34] = 32147
          "0111110010100011" when "100011", -- t[35] = 31907
          "0111101110110110" when "100100", -- t[36] = 31670
          "0111101011001111" when "100101", -- t[37] = 31439
          "0111100111101100" when "100110", -- t[38] = 31212
          "0111100100001101" when "100111", -- t[39] = 30989
          "0111100000110010" when "101000", -- t[40] = 30770
          "0111011101011100" when "101001", -- t[41] = 30556
          "0111011010001001" when "101010", -- t[42] = 30345
          "0111010110111010" when "101011", -- t[43] = 30138
          "0111010011101111" when "101100", -- t[44] = 29935
          "0111010000100111" when "101101", -- t[45] = 29735
          "0111001101100011" when "101110", -- t[46] = 29539
          "0111001010100010" when "101111", -- t[47] = 29346
          "0111000111100100" when "110000", -- t[48] = 29156
          "0111000100101010" when "110001", -- t[49] = 28970
          "0111000001110010" when "110010", -- t[50] = 28786
          "0110111110111110" when "110011", -- t[51] = 28606
          "0110111100001101" when "110100", -- t[52] = 28429
          "0110111001011110" when "110101", -- t[53] = 28254
          "0110110110110010" when "110110", -- t[54] = 28082
          "0110110100001001" when "110111", -- t[55] = 27913
          "0110110001100010" when "111000", -- t[56] = 27746
          "0110101110111110" when "111001", -- t[57] = 27582
          "0110101100011101" when "111010", -- t[58] = 27421
          "0110101001111110" when "111011", -- t[59] = 27262
          "0110100111100001" when "111100", -- t[60] = 27105
          "0110100101000111" when "111101", -- t[61] = 26951
          "0110100010101111" when "111110", -- t[62] = 26799
          "0110100000011001" when "111111", -- t[63] = 26649
          "----------------" when others;

  r(15 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 6; mu_1 = 6; lambda_1 = 6.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_12_t1_pow is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_log_log_12_t1_pow is
  signal pp0 : std_logic_vector(4 downto 0);
  signal r0 : std_logic_vector(4 downto 0);
begin
  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(4 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 6; wO_1,1 = 10.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_12_t1_t1 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of fp_log_log_12_t1_t1 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a;

  with x select
    r <= "1001101001" when "000000", -- t[0] = 617
         "1001010001" when "000001", -- t[1] = 593
         "1000111100" when "000010", -- t[2] = 572
         "1000100111" when "000011", -- t[3] = 551
         "1000010100" when "000100", -- t[4] = 532
         "1000000010" when "000101", -- t[5] = 514
         "0111110001" when "000110", -- t[6] = 497
         "0111100001" when "000111", -- t[7] = 481
         "0111010010" when "001000", -- t[8] = 466
         "0111000100" when "001001", -- t[9] = 452
         "0110110110" when "001010", -- t[10] = 438
         "0110101001" when "001011", -- t[11] = 425
         "0110011101" when "001100", -- t[12] = 413
         "0110010001" when "001101", -- t[13] = 401
         "0110000110" when "001110", -- t[14] = 390
         "0101111011" when "001111", -- t[15] = 379
         "0101110001" when "010000", -- t[16] = 369
         "0101100111" when "010001", -- t[17] = 359
         "0101011110" when "010010", -- t[18] = 350
         "0101010101" when "010011", -- t[19] = 341
         "0101001101" when "010100", -- t[20] = 333
         "0101000101" when "010101", -- t[21] = 325
         "0100111101" when "010110", -- t[22] = 317
         "0100110101" when "010111", -- t[23] = 309
         "0100101110" when "011000", -- t[24] = 302
         "0100100111" when "011001", -- t[25] = 295
         "0100100001" when "011010", -- t[26] = 289
         "0100011010" when "011011", -- t[27] = 282
         "0100010100" when "011100", -- t[28] = 276
         "0100001110" when "011101", -- t[29] = 270
         "0100001000" when "011110", -- t[30] = 264
         "0100000011" when "011111", -- t[31] = 259
         "0011111101" when "100000", -- t[32] = 253
         "0011111000" when "100001", -- t[33] = 248
         "0011110011" when "100010", -- t[34] = 243
         "0011101110" when "100011", -- t[35] = 238
         "0011101010" when "100100", -- t[36] = 234
         "0011100101" when "100101", -- t[37] = 229
         "0011100001" when "100110", -- t[38] = 225
         "0011011101" when "100111", -- t[39] = 221
         "0011011001" when "101000", -- t[40] = 217
         "0011010101" when "101001", -- t[41] = 213
         "0011010001" when "101010", -- t[42] = 209
         "0011001101" when "101011", -- t[43] = 205
         "0011001001" when "101100", -- t[44] = 201
         "0011000110" when "101101", -- t[45] = 198
         "0011000011" when "101110", -- t[46] = 195
         "0010111111" when "101111", -- t[47] = 191
         "0010111100" when "110000", -- t[48] = 188
         "0010111001" when "110001", -- t[49] = 185
         "0010110110" when "110010", -- t[50] = 182
         "0010110011" when "110011", -- t[51] = 179
         "0010110000" when "110100", -- t[52] = 176
         "0010101101" when "110101", -- t[53] = 173
         "0010101010" when "110110", -- t[54] = 170
         "0010101000" when "110111", -- t[55] = 168
         "0010100101" when "111000", -- t[56] = 165
         "0010100011" when "111001", -- t[57] = 163
         "0010100000" when "111010", -- t[58] = 160
         "0010011110" when "111011", -- t[59] = 158
         "0010011011" when "111100", -- t[60] = 155
         "0010011001" when "111101", -- t[61] = 153
         "0010010111" when "111110", -- t[62] = 151
         "0010010101" when "111111", -- t[63] = 149
         "----------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_2.
-- Decomposition:
--   alpha_1,2 = 4; sigma'_1,2 = 1; wO_1,2 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_12_t1_t2 is
  port ( a : in  std_logic_vector(3 downto 0);
         s : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_log_log_12_t1_t2 is
  signal x : std_logic_vector(4 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0100" when "00000", -- t[0] = 4
         "1101" when "00001", -- t[1] = 13
         "0011" when "00010", -- t[2] = 3
         "1011" when "00011", -- t[3] = 11
         "0011" when "00100", -- t[4] = 3
         "1010" when "00101", -- t[5] = 10
         "0011" when "00110", -- t[6] = 3
         "1001" when "00111", -- t[7] = 9
         "0010" when "01000", -- t[8] = 2
         "1000" when "01001", -- t[9] = 8
         "0010" when "01010", -- t[10] = 2
         "0111" when "01011", -- t[11] = 7
         "0010" when "01100", -- t[12] = 2
         "0110" when "01101", -- t[13] = 6
         "0010" when "01110", -- t[14] = 2
         "0110" when "01111", -- t[15] = 6
         "0001" when "10000", -- t[16] = 1
         "0101" when "10001", -- t[17] = 5
         "0001" when "10010", -- t[18] = 1
         "0101" when "10011", -- t[19] = 5
         "0001" when "10100", -- t[20] = 1
         "0100" when "10101", -- t[21] = 4
         "0001" when "10110", -- t[22] = 1
         "0100" when "10111", -- t[23] = 4
         "0001" when "11000", -- t[24] = 1
         "0100" when "11001", -- t[25] = 4
         "0001" when "11010", -- t[26] = 1
         "0100" when "11011", -- t[27] = 4
         "0001" when "11100", -- t[28] = 1
         "0011" when "11101", -- t[29] = 3
         "0001" when "11110", -- t[30] = 1
         "0011" when "11111", -- t[31] = 3
         "----" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 6; beta_1 = 6; lambda_1 = 6;  m_1 = 2;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 6; rho_1,1 = 0; sigma_1,1 = 4; wO_1,1 = 10;
--   Q_1,2 (ROM):  alpha_1,2 = 4; rho_1,2 = 4; sigma_1,2 = 2; wO_1,2 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_12_t1 is
  port ( a : in  std_logic_vector(5 downto 0);
         b : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of fp_log_log_12_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(4 downto 0);
  signal s      : std_logic_vector(5 downto 0);
  component fp_log_log_12_t1_pow is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  signal a_1    : std_logic_vector(5 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(2 downto 0);
  signal k_1    : std_logic_vector(9 downto 0);
  signal r0_1   : std_logic_vector(14 downto 0);
  signal r_1    : std_logic_vector(15 downto 0);
  component fp_log_log_12_t1_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  signal a_2    : std_logic_vector(3 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(0 downto 0);
  signal r0_2   : std_logic_vector(3 downto 0);
  signal r_2    : std_logic_vector(15 downto 0);
  component fp_log_log_12_t1_t2 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;
begin
  sign <= not b(5);
  b0 <= b(4 downto 0) xor (4 downto 0 => sign);

  pow : fp_log_log_12_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(5 downto 0);
  sign_1 <= not s(5);
  s_1 <= s(4 downto 2) xor (4 downto 2 => sign_1);
  t_1 : fp_log_log_12_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(9 downto 0) <=
    r0_1(14 downto 5) xor (14 downto 5 => (not (sign xor sign_1)));
  r_1(15 downto 10) <= (15 downto 10 => (not (sign xor sign_1)));

  a_2 <= a(5 downto 2);
  sign_2 <= not s(1);
  s_2 <= s(0 downto 0) xor (0 downto 0 => sign_2);
  t_2 : fp_log_log_12_t1_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(3 downto 0) <=
    r0_2 xor (3 downto 0 => (not (sign xor sign_2)));
  r_2(15 downto 4) <= (15 downto 4 => (not (sign xor sign_2)));

  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_12 is
  port ( x : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of fp_log_log_12 is
  signal a_0 : std_logic_vector(5 downto 0);
  signal r_0 : std_logic_vector(15 downto 0);
  component fp_log_log_12_t0 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(15 downto 0) );
  end component;

  signal a_1 : std_logic_vector(5 downto 0);
  signal b_1 : std_logic_vector(5 downto 0);
  signal r_1 : std_logic_vector(15 downto 0);
  component fp_log_log_12_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           b : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(15 downto 0) );
  end component;

begin
  a_0 <= x(11 downto 6);
  t_0 : fp_log_log_12_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(11 downto 6);
  b_1 <= x(5 downto 0);
  t_1 : fp_log_log_12_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  r <= r_0 + r_1;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 13; wO = 13.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 6;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 7; beta_1 = 6.
-- Guard bits: g = 3.
-- Command line: logfp 13 13 1   rom 7 0   pm 7 6  ah 6 6 6  1 1  7 4 0  3 2 4


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 17.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_13_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of fp_log_log_13_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(16 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110000110110010" when "0000000", -- t[0] = 90546
          "10101111101001010" when "0000001", -- t[1] = 89930
          "10101110011101101" when "0000010", -- t[2] = 89325
          "10101101010011100" when "0000011", -- t[3] = 88732
          "10101100001010101" when "0000100", -- t[4] = 88149
          "10101011000011010" when "0000101", -- t[5] = 87578
          "10101001111101001" when "0000110", -- t[6] = 87017
          "10101000111000001" when "0000111", -- t[7] = 86465
          "10100111110100100" when "0001000", -- t[8] = 85924
          "10100110110010000" when "0001001", -- t[9] = 85392
          "10100101110000101" when "0001010", -- t[10] = 84869
          "10100100110000011" when "0001011", -- t[11] = 84355
          "10100011110001001" when "0001100", -- t[12] = 83849
          "10100010110011000" when "0001101", -- t[13] = 83352
          "10100001110101111" when "0001110", -- t[14] = 82863
          "10100000111001110" when "0001111", -- t[15] = 82382
          "10011111111110101" when "0010000", -- t[16] = 81909
          "10011111000100011" when "0010001", -- t[17] = 81443
          "10011110001011000" when "0010010", -- t[18] = 80984
          "10011101010010100" when "0010011", -- t[19] = 80532
          "10011100011011000" when "0010100", -- t[20] = 80088
          "10011011100100010" when "0010101", -- t[21] = 79650
          "10011010101110011" when "0010110", -- t[22] = 79219
          "10011001111001010" when "0010111", -- t[23] = 78794
          "10011001000100111" when "0011000", -- t[24] = 78375
          "10011000010001010" when "0011001", -- t[25] = 77962
          "10010111011110100" when "0011010", -- t[26] = 77556
          "10010110101100011" when "0011011", -- t[27] = 77155
          "10010101111010111" when "0011100", -- t[28] = 76759
          "10010101001010010" when "0011101", -- t[29] = 76370
          "10010100011010001" when "0011110", -- t[30] = 75985
          "10010011101010110" when "0011111", -- t[31] = 75606
          "10010010111100000" when "0100000", -- t[32] = 75232
          "10010010001101111" when "0100001", -- t[33] = 74863
          "10010001100000011" when "0100010", -- t[34] = 74499
          "10010000110011100" when "0100011", -- t[35] = 74140
          "10010000000111001" when "0100100", -- t[36] = 73785
          "10001111011011011" when "0100101", -- t[37] = 73435
          "10001110110000001" when "0100110", -- t[38] = 73089
          "10001110000101100" when "0100111", -- t[39] = 72748
          "10001101011011011" when "0101000", -- t[40] = 72411
          "10001100110001110" when "0101001", -- t[41] = 72078
          "10001100001000110" when "0101010", -- t[42] = 71750
          "10001011100000001" when "0101011", -- t[43] = 71425
          "10001010111000001" when "0101100", -- t[44] = 71105
          "10001010010000100" when "0101101", -- t[45] = 70788
          "10001001101001011" when "0101110", -- t[46] = 70475
          "10001001000010110" when "0101111", -- t[47] = 70166
          "10001000011100100" when "0110000", -- t[48] = 69860
          "10000111110110110" when "0110001", -- t[49] = 69558
          "10000111010001100" when "0110010", -- t[50] = 69260
          "10000110101100100" when "0110011", -- t[51] = 68964
          "10000110001000001" when "0110100", -- t[52] = 68673
          "10000101100100000" when "0110101", -- t[53] = 68384
          "10000101000000011" when "0110110", -- t[54] = 68099
          "10000100011101001" when "0110111", -- t[55] = 67817
          "10000011111010010" when "0111000", -- t[56] = 67538
          "10000011010111110" when "0111001", -- t[57] = 67262
          "10000010110101101" when "0111010", -- t[58] = 66989
          "10000010010011111" when "0111011", -- t[59] = 66719
          "10000001110010100" when "0111100", -- t[60] = 66452
          "10000001010001100" when "0111101", -- t[61] = 66188
          "10000000110000110" when "0111110", -- t[62] = 65926
          "10000000010000100" when "0111111", -- t[63] = 65668
          "01111111110000011" when "1000000", -- t[64] = 65411
          "01111111010000110" when "1000001", -- t[65] = 65158
          "01111110110001011" when "1000010", -- t[66] = 64907
          "01111110010010011" when "1000011", -- t[67] = 64659
          "01111101110011101" when "1000100", -- t[68] = 64413
          "01111101010101010" when "1000101", -- t[69] = 64170
          "01111100110111001" when "1000110", -- t[70] = 63929
          "01111100011001011" when "1000111", -- t[71] = 63691
          "01111011111011111" when "1001000", -- t[72] = 63455
          "01111011011110101" when "1001001", -- t[73] = 63221
          "01111011000001101" when "1001010", -- t[74] = 62989
          "01111010100101000" when "1001011", -- t[75] = 62760
          "01111010001000101" when "1001100", -- t[76] = 62533
          "01111001101100100" when "1001101", -- t[77] = 62308
          "01111001010000101" when "1001110", -- t[78] = 62085
          "01111000110101001" when "1001111", -- t[79] = 61865
          "01111000011001110" when "1010000", -- t[80] = 61646
          "01110111111110101" when "1010001", -- t[81] = 61429
          "01110111100011111" when "1010010", -- t[82] = 61215
          "01110111001001010" when "1010011", -- t[83] = 61002
          "01110110101110111" when "1010100", -- t[84] = 60791
          "01110110010100111" when "1010101", -- t[85] = 60583
          "01110101111011000" when "1010110", -- t[86] = 60376
          "01110101100001011" when "1010111", -- t[87] = 60171
          "01110101000111111" when "1011000", -- t[88] = 59967
          "01110100101110110" when "1011001", -- t[89] = 59766
          "01110100010101110" when "1011010", -- t[90] = 59566
          "01110011111101000" when "1011011", -- t[91] = 59368
          "01110011100100100" when "1011100", -- t[92] = 59172
          "01110011001100001" when "1011101", -- t[93] = 58977
          "01110010110100001" when "1011110", -- t[94] = 58785
          "01110010011100001" when "1011111", -- t[95] = 58593
          "01110010000100100" when "1100000", -- t[96] = 58404
          "01110001101101000" when "1100001", -- t[97] = 58216
          "01110001010101101" when "1100010", -- t[98] = 58029
          "01110000111110100" when "1100011", -- t[99] = 57844
          "01110000100111101" when "1100100", -- t[100] = 57661
          "01110000010000111" when "1100101", -- t[101] = 57479
          "01101111111010011" when "1100110", -- t[102] = 57299
          "01101111100100000" when "1100111", -- t[103] = 57120
          "01101111001101111" when "1101000", -- t[104] = 56943
          "01101110110111111" when "1101001", -- t[105] = 56767
          "01101110100010000" when "1101010", -- t[106] = 56592
          "01101110001100011" when "1101011", -- t[107] = 56419
          "01101101110110111" when "1101100", -- t[108] = 56247
          "01101101100001101" when "1101101", -- t[109] = 56077
          "01101101001100011" when "1101110", -- t[110] = 55907
          "01101100110111100" when "1101111", -- t[111] = 55740
          "01101100100010101" when "1110000", -- t[112] = 55573
          "01101100001110000" when "1110001", -- t[113] = 55408
          "01101011111001100" when "1110010", -- t[114] = 55244
          "01101011100101001" when "1110011", -- t[115] = 55081
          "01101011010001000" when "1110100", -- t[116] = 54920
          "01101010111101000" when "1110101", -- t[117] = 54760
          "01101010101001001" when "1110110", -- t[118] = 54601
          "01101010010101011" when "1110111", -- t[119] = 54443
          "01101010000001110" when "1111000", -- t[120] = 54286
          "01101001101110011" when "1111001", -- t[121] = 54131
          "01101001011011000" when "1111010", -- t[122] = 53976
          "01101001000111111" when "1111011", -- t[123] = 53823
          "01101000110100111" when "1111100", -- t[124] = 53671
          "01101000100010000" when "1111101", -- t[125] = 53520
          "01101000001111010" when "1111110", -- t[126] = 53370
          "01100111111100101" when "1111111", -- t[127] = 53221
          "-----------------" when others;

  r(16 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 6; mu_1 = 6; lambda_1 = 6.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_13_t1_pow is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_log_log_13_t1_pow is
  signal pp0 : std_logic_vector(4 downto 0);
  signal r0 : std_logic_vector(4 downto 0);
begin
  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(4 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 7; wO_1,1 = 10.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_13_t1_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of fp_log_log_13_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "1001101110" when "0000000", -- t[0] = 622
         "1001100010" when "0000001", -- t[1] = 610
         "1001010111" when "0000010", -- t[2] = 599
         "1001001100" when "0000011", -- t[3] = 588
         "1001000001" when "0000100", -- t[4] = 577
         "1000110110" when "0000101", -- t[5] = 566
         "1000101100" when "0000110", -- t[6] = 556
         "1000100010" when "0000111", -- t[7] = 546
         "1000011001" when "0001000", -- t[8] = 537
         "1000010000" when "0001001", -- t[9] = 528
         "1000000111" when "0001010", -- t[10] = 519
         "0111111110" when "0001011", -- t[11] = 510
         "0111110101" when "0001100", -- t[12] = 501
         "0111101101" when "0001101", -- t[13] = 493
         "0111100101" when "0001110", -- t[14] = 485
         "0111011101" when "0001111", -- t[15] = 477
         "0111010110" when "0010000", -- t[16] = 470
         "0111001110" when "0010001", -- t[17] = 462
         "0111000111" when "0010010", -- t[18] = 455
         "0111000000" when "0010011", -- t[19] = 448
         "0110111001" when "0010100", -- t[20] = 441
         "0110110011" when "0010101", -- t[21] = 435
         "0110101100" when "0010110", -- t[22] = 428
         "0110100110" when "0010111", -- t[23] = 422
         "0110100000" when "0011000", -- t[24] = 416
         "0110011010" when "0011001", -- t[25] = 410
         "0110010100" when "0011010", -- t[26] = 404
         "0110001110" when "0011011", -- t[27] = 398
         "0110001001" when "0011100", -- t[28] = 393
         "0110000011" when "0011101", -- t[29] = 387
         "0101111110" when "0011110", -- t[30] = 382
         "0101111001" when "0011111", -- t[31] = 377
         "0101110011" when "0100000", -- t[32] = 371
         "0101101111" when "0100001", -- t[33] = 367
         "0101101010" when "0100010", -- t[34] = 362
         "0101100101" when "0100011", -- t[35] = 357
         "0101100000" when "0100100", -- t[36] = 352
         "0101011100" when "0100101", -- t[37] = 348
         "0101010111" when "0100110", -- t[38] = 343
         "0101010011" when "0100111", -- t[39] = 339
         "0101001111" when "0101000", -- t[40] = 335
         "0101001011" when "0101001", -- t[41] = 331
         "0101000111" when "0101010", -- t[42] = 327
         "0101000011" when "0101011", -- t[43] = 323
         "0100111111" when "0101100", -- t[44] = 319
         "0100111011" when "0101101", -- t[45] = 315
         "0100110111" when "0101110", -- t[46] = 311
         "0100110011" when "0101111", -- t[47] = 307
         "0100110000" when "0110000", -- t[48] = 304
         "0100101100" when "0110001", -- t[49] = 300
         "0100101001" when "0110010", -- t[50] = 297
         "0100100101" when "0110011", -- t[51] = 293
         "0100100010" when "0110100", -- t[52] = 290
         "0100011111" when "0110101", -- t[53] = 287
         "0100011100" when "0110110", -- t[54] = 284
         "0100011001" when "0110111", -- t[55] = 281
         "0100010101" when "0111000", -- t[56] = 277
         "0100010010" when "0111001", -- t[57] = 274
         "0100001111" when "0111010", -- t[58] = 271
         "0100001101" when "0111011", -- t[59] = 269
         "0100001010" when "0111100", -- t[60] = 266
         "0100000111" when "0111101", -- t[61] = 263
         "0100000100" when "0111110", -- t[62] = 260
         "0100000001" when "0111111", -- t[63] = 257
         "0011111111" when "1000000", -- t[64] = 255
         "0011111100" when "1000001", -- t[65] = 252
         "0011111001" when "1000010", -- t[66] = 249
         "0011110111" when "1000011", -- t[67] = 247
         "0011110100" when "1000100", -- t[68] = 244
         "0011110010" when "1000101", -- t[69] = 242
         "0011110000" when "1000110", -- t[70] = 240
         "0011101101" when "1000111", -- t[71] = 237
         "0011101011" when "1001000", -- t[72] = 235
         "0011101001" when "1001001", -- t[73] = 233
         "0011100110" when "1001010", -- t[74] = 230
         "0011100100" when "1001011", -- t[75] = 228
         "0011100010" when "1001100", -- t[76] = 226
         "0011100000" when "1001101", -- t[77] = 224
         "0011011110" when "1001110", -- t[78] = 222
         "0011011100" when "1001111", -- t[79] = 220
         "0011011010" when "1010000", -- t[80] = 218
         "0011011000" when "1010001", -- t[81] = 216
         "0011010110" when "1010010", -- t[82] = 214
         "0011010100" when "1010011", -- t[83] = 212
         "0011010010" when "1010100", -- t[84] = 210
         "0011010000" when "1010101", -- t[85] = 208
         "0011001110" when "1010110", -- t[86] = 206
         "0011001100" when "1010111", -- t[87] = 204
         "0011001010" when "1011000", -- t[88] = 202
         "0011001001" when "1011001", -- t[89] = 201
         "0011000111" when "1011010", -- t[90] = 199
         "0011000101" when "1011011", -- t[91] = 197
         "0011000011" when "1011100", -- t[92] = 195
         "0011000010" when "1011101", -- t[93] = 194
         "0011000000" when "1011110", -- t[94] = 192
         "0010111110" when "1011111", -- t[95] = 190
         "0010111101" when "1100000", -- t[96] = 189
         "0010111011" when "1100001", -- t[97] = 187
         "0010111010" when "1100010", -- t[98] = 186
         "0010111000" when "1100011", -- t[99] = 184
         "0010110111" when "1100100", -- t[100] = 183
         "0010110101" when "1100101", -- t[101] = 181
         "0010110100" when "1100110", -- t[102] = 180
         "0010110010" when "1100111", -- t[103] = 178
         "0010110001" when "1101000", -- t[104] = 177
         "0010101111" when "1101001", -- t[105] = 175
         "0010101110" when "1101010", -- t[106] = 174
         "0010101100" when "1101011", -- t[107] = 172
         "0010101011" when "1101100", -- t[108] = 171
         "0010101010" when "1101101", -- t[109] = 170
         "0010101000" when "1101110", -- t[110] = 168
         "0010100111" when "1101111", -- t[111] = 167
         "0010100110" when "1110000", -- t[112] = 166
         "0010100101" when "1110001", -- t[113] = 165
         "0010100011" when "1110010", -- t[114] = 163
         "0010100010" when "1110011", -- t[115] = 162
         "0010100001" when "1110100", -- t[116] = 161
         "0010100000" when "1110101", -- t[117] = 160
         "0010011110" when "1110110", -- t[118] = 158
         "0010011101" when "1110111", -- t[119] = 157
         "0010011100" when "1111000", -- t[120] = 156
         "0010011011" when "1111001", -- t[121] = 155
         "0010011010" when "1111010", -- t[122] = 154
         "0010011001" when "1111011", -- t[123] = 153
         "0010011000" when "1111100", -- t[124] = 152
         "0010010110" when "1111101", -- t[125] = 150
         "0010010101" when "1111110", -- t[126] = 149
         "0010010100" when "1111111", -- t[127] = 148
         "----------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_2.
-- Decomposition:
--   alpha_1,2 = 3; sigma'_1,2 = 1; wO_1,2 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_13_t1_t2 is
  port ( a : in  std_logic_vector(2 downto 0);
         s : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of fp_log_log_13_t1_t2 is
  signal x : std_logic_vector(3 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0100" when "0000", -- t[0] = 4
         "1100" when "0001", -- t[1] = 12
         "0011" when "0010", -- t[2] = 3
         "1001" when "0011", -- t[3] = 9
         "0010" when "0100", -- t[4] = 2
         "0111" when "0101", -- t[5] = 7
         "0010" when "0110", -- t[6] = 2
         "0110" when "0111", -- t[7] = 6
         "0001" when "1000", -- t[8] = 1
         "0101" when "1001", -- t[9] = 5
         "0001" when "1010", -- t[10] = 1
         "0100" when "1011", -- t[11] = 4
         "0001" when "1100", -- t[12] = 1
         "0100" when "1101", -- t[13] = 4
         "0001" when "1110", -- t[14] = 1
         "0011" when "1111", -- t[15] = 3
         "----" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 7; beta_1 = 6; lambda_1 = 6;  m_1 = 2;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 7; rho_1,1 = 0; sigma_1,1 = 4; wO_1,1 = 10;
--   Q_1,2 (ROM):  alpha_1,2 = 3; rho_1,2 = 4; sigma_1,2 = 2; wO_1,2 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_13_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of fp_log_log_13_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(4 downto 0);
  signal s      : std_logic_vector(5 downto 0);
  component fp_log_log_13_t1_pow is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(2 downto 0);
  signal k_1    : std_logic_vector(9 downto 0);
  signal r0_1   : std_logic_vector(14 downto 0);
  signal r_1    : std_logic_vector(16 downto 0);
  component fp_log_log_13_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  signal a_2    : std_logic_vector(2 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(0 downto 0);
  signal r0_2   : std_logic_vector(3 downto 0);
  signal r_2    : std_logic_vector(16 downto 0);
  component fp_log_log_13_t1_t2 is
    port ( a : in  std_logic_vector(2 downto 0);
           s : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;
begin
  sign <= not b(5);
  b0 <= b(4 downto 0) xor (4 downto 0 => sign);

  pow : fp_log_log_13_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(5);
  s_1 <= s(4 downto 2) xor (4 downto 2 => sign_1);
  t_1 : fp_log_log_13_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(9 downto 0) <=
    r0_1(14 downto 5) xor (14 downto 5 => (not (sign xor sign_1)));
  r_1(16 downto 10) <= (16 downto 10 => (not (sign xor sign_1)));

  a_2 <= a(6 downto 4);
  sign_2 <= not s(1);
  s_2 <= s(0 downto 0) xor (0 downto 0 => sign_2);
  t_2 : fp_log_log_13_t1_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(3 downto 0) <=
    r0_2 xor (3 downto 0 => (not (sign xor sign_2)));
  r_2(16 downto 4) <= (16 downto 4 => (not (sign xor sign_2)));

  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_13 is
  port ( x : in  std_logic_vector(12 downto 0);
         r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of fp_log_log_13 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(16 downto 0);
  component fp_log_log_13_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(16 downto 0) );
  end component;

  signal a_1 : std_logic_vector(6 downto 0);
  signal b_1 : std_logic_vector(5 downto 0);
  signal r_1 : std_logic_vector(16 downto 0);
  component fp_log_log_13_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(16 downto 0) );
  end component;

begin
  a_0 <= x(12 downto 6);
  t_0 : fp_log_log_13_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(12 downto 6);
  b_1 <= x(5 downto 0);
  t_1 : fp_log_log_13_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  r <= r_0 + r_1;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 14; wO = 14.
-- Order-1 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 7;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 7; beta_1 = 7.
-- Guard bits: g = 2.
-- Command line: logfp 14 14 1   rom 7 0   pm 7 7  ah 7 7 7  1 0  7 7 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 17.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_14_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of fp_log_log_14_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(16 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110000110101111" when "0000000", -- t[0] = 90543
          "10101111101000111" when "0000001", -- t[1] = 89927
          "10101110011101010" when "0000010", -- t[2] = 89322
          "10101101010011001" when "0000011", -- t[3] = 88729
          "10101100001010011" when "0000100", -- t[4] = 88147
          "10101011000010111" when "0000101", -- t[5] = 87575
          "10101001111100110" when "0000110", -- t[6] = 87014
          "10101000110111111" when "0000111", -- t[7] = 86463
          "10100111110100001" when "0001000", -- t[8] = 85921
          "10100110110001101" when "0001001", -- t[9] = 85389
          "10100101110000010" when "0001010", -- t[10] = 84866
          "10100100110000000" when "0001011", -- t[11] = 84352
          "10100011110000111" when "0001100", -- t[12] = 83847
          "10100010110010110" when "0001101", -- t[13] = 83350
          "10100001110101101" when "0001110", -- t[14] = 82861
          "10100000111001100" when "0001111", -- t[15] = 82380
          "10011111111110010" when "0010000", -- t[16] = 81906
          "10011111000100000" when "0010001", -- t[17] = 81440
          "10011110001010110" when "0010010", -- t[18] = 80982
          "10011101010010010" when "0010011", -- t[19] = 80530
          "10011100011010110" when "0010100", -- t[20] = 80086
          "10011011100100000" when "0010101", -- t[21] = 79648
          "10011010101110000" when "0010110", -- t[22] = 79216
          "10011001111001000" when "0010111", -- t[23] = 78792
          "10011001000100101" when "0011000", -- t[24] = 78373
          "10011000010001000" when "0011001", -- t[25] = 77960
          "10010111011110010" when "0011010", -- t[26] = 77554
          "10010110101100001" when "0011011", -- t[27] = 77153
          "10010101111010101" when "0011100", -- t[28] = 76757
          "10010101001010000" when "0011101", -- t[29] = 76368
          "10010100011001111" when "0011110", -- t[30] = 75983
          "10010011101010100" when "0011111", -- t[31] = 75604
          "10010010111011110" when "0100000", -- t[32] = 75230
          "10010010001101101" when "0100001", -- t[33] = 74861
          "10010001100000001" when "0100010", -- t[34] = 74497
          "10010000110011010" when "0100011", -- t[35] = 74138
          "10010000000110111" when "0100100", -- t[36] = 73783
          "10001111011011001" when "0100101", -- t[37] = 73433
          "10001110101111111" when "0100110", -- t[38] = 73087
          "10001110000101010" when "0100111", -- t[39] = 72746
          "10001101011011001" when "0101000", -- t[40] = 72409
          "10001100110001101" when "0101001", -- t[41] = 72077
          "10001100001000100" when "0101010", -- t[42] = 71748
          "10001011100000000" when "0101011", -- t[43] = 71424
          "10001010110111111" when "0101100", -- t[44] = 71103
          "10001010010000010" when "0101101", -- t[45] = 70786
          "10001001101001001" when "0101110", -- t[46] = 70473
          "10001001000010100" when "0101111", -- t[47] = 70164
          "10001000011100010" when "0110000", -- t[48] = 69858
          "10000111110110100" when "0110001", -- t[49] = 69556
          "10000111010001010" when "0110010", -- t[50] = 69258
          "10000110101100011" when "0110011", -- t[51] = 68963
          "10000110000111111" when "0110100", -- t[52] = 68671
          "10000101100011111" when "0110101", -- t[53] = 68383
          "10000101000000001" when "0110110", -- t[54] = 68097
          "10000100011100111" when "0110111", -- t[55] = 67815
          "10000011111010000" when "0111000", -- t[56] = 67536
          "10000011010111100" when "0111001", -- t[57] = 67260
          "10000010110101011" when "0111010", -- t[58] = 66987
          "10000010010011101" when "0111011", -- t[59] = 66717
          "10000001110010010" when "0111100", -- t[60] = 66450
          "10000001010001010" when "0111101", -- t[61] = 66186
          "10000000110000101" when "0111110", -- t[62] = 65925
          "10000000010000010" when "0111111", -- t[63] = 65666
          "01111111110000010" when "1000000", -- t[64] = 65410
          "01111111010000101" when "1000001", -- t[65] = 65157
          "01111110110001010" when "1000010", -- t[66] = 64906
          "01111110010010010" when "1000011", -- t[67] = 64658
          "01111101110011100" when "1000100", -- t[68] = 64412
          "01111101010101001" when "1000101", -- t[69] = 64169
          "01111100110111000" when "1000110", -- t[70] = 63928
          "01111100011001001" when "1000111", -- t[71] = 63689
          "01111011111011101" when "1001000", -- t[72] = 63453
          "01111011011110100" when "1001001", -- t[73] = 63220
          "01111011000001100" when "1001010", -- t[74] = 62988
          "01111010100100111" when "1001011", -- t[75] = 62759
          "01111010001000100" when "1001100", -- t[76] = 62532
          "01111001101100011" when "1001101", -- t[77] = 62307
          "01111001010000100" when "1001110", -- t[78] = 62084
          "01111000110100111" when "1001111", -- t[79] = 61863
          "01111000011001101" when "1010000", -- t[80] = 61645
          "01110111111110100" when "1010001", -- t[81] = 61428
          "01110111100011101" when "1010010", -- t[82] = 61213
          "01110111001001001" when "1010011", -- t[83] = 61001
          "01110110101110110" when "1010100", -- t[84] = 60790
          "01110110010100101" when "1010101", -- t[85] = 60581
          "01110101111010110" when "1010110", -- t[86] = 60374
          "01110101100001001" when "1010111", -- t[87] = 60169
          "01110101000111110" when "1011000", -- t[88] = 59966
          "01110100101110101" when "1011001", -- t[89] = 59765
          "01110100010101101" when "1011010", -- t[90] = 59565
          "01110011111100111" when "1011011", -- t[91] = 59367
          "01110011100100011" when "1011100", -- t[92] = 59171
          "01110011001100000" when "1011101", -- t[93] = 58976
          "01110010110011111" when "1011110", -- t[94] = 58783
          "01110010011100000" when "1011111", -- t[95] = 58592
          "01110010000100010" when "1100000", -- t[96] = 58402
          "01110001101100110" when "1100001", -- t[97] = 58214
          "01110001010101100" when "1100010", -- t[98] = 58028
          "01110000111110011" when "1100011", -- t[99] = 57843
          "01110000100111100" when "1100100", -- t[100] = 57660
          "01110000010000110" when "1100101", -- t[101] = 57478
          "01101111111010010" when "1100110", -- t[102] = 57298
          "01101111100011111" when "1100111", -- t[103] = 57119
          "01101111001101101" when "1101000", -- t[104] = 56941
          "01101110110111101" when "1101001", -- t[105] = 56765
          "01101110100001111" when "1101010", -- t[106] = 56591
          "01101110001100010" when "1101011", -- t[107] = 56418
          "01101101110110110" when "1101100", -- t[108] = 56246
          "01101101100001011" when "1101101", -- t[109] = 56075
          "01101101001100010" when "1101110", -- t[110] = 55906
          "01101100110111010" when "1101111", -- t[111] = 55738
          "01101100100010100" when "1110000", -- t[112] = 55572
          "01101100001101111" when "1110001", -- t[113] = 55407
          "01101011111001011" when "1110010", -- t[114] = 55243
          "01101011100101000" when "1110011", -- t[115] = 55080
          "01101011010000111" when "1110100", -- t[116] = 54919
          "01101010111100110" when "1110101", -- t[117] = 54758
          "01101010101000111" when "1110110", -- t[118] = 54599
          "01101010010101010" when "1110111", -- t[119] = 54442
          "01101010000001101" when "1111000", -- t[120] = 54285
          "01101001101110010" when "1111001", -- t[121] = 54130
          "01101001011010111" when "1111010", -- t[122] = 53975
          "01101001000111110" when "1111011", -- t[123] = 53822
          "01101000110100110" when "1111100", -- t[124] = 53670
          "01101000100001111" when "1111101", -- t[125] = 53519
          "01101000001111001" when "1111110", -- t[126] = 53369
          "01100111111100100" when "1111111", -- t[127] = 53220
          "-----------------" when others;

  r(16 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 7; mu_1 = 7; lambda_1 = 7.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_14_t1_pow is
  port ( x : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_log_log_14_t1_pow is
  signal pp0 : std_logic_vector(5 downto 0);
  signal r0 : std_logic_vector(5 downto 0);
begin
  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(5 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 7; wO_1,1 = 10.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_14_t1_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of fp_log_log_14_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "1001101110" when "0000000", -- t[0] = 622
         "1001100010" when "0000001", -- t[1] = 610
         "1001010111" when "0000010", -- t[2] = 599
         "1001001100" when "0000011", -- t[3] = 588
         "1001000001" when "0000100", -- t[4] = 577
         "1000110110" when "0000101", -- t[5] = 566
         "1000101100" when "0000110", -- t[6] = 556
         "1000100010" when "0000111", -- t[7] = 546
         "1000011001" when "0001000", -- t[8] = 537
         "1000001111" when "0001001", -- t[9] = 527
         "1000000110" when "0001010", -- t[10] = 518
         "0111111110" when "0001011", -- t[11] = 510
         "0111110101" when "0001100", -- t[12] = 501
         "0111101101" when "0001101", -- t[13] = 493
         "0111100101" when "0001110", -- t[14] = 485
         "0111011101" when "0001111", -- t[15] = 477
         "0111010110" when "0010000", -- t[16] = 470
         "0111001110" when "0010001", -- t[17] = 462
         "0111000111" when "0010010", -- t[18] = 455
         "0111000000" when "0010011", -- t[19] = 448
         "0110111001" when "0010100", -- t[20] = 441
         "0110110011" when "0010101", -- t[21] = 435
         "0110101100" when "0010110", -- t[22] = 428
         "0110100110" when "0010111", -- t[23] = 422
         "0110100000" when "0011000", -- t[24] = 416
         "0110011010" when "0011001", -- t[25] = 410
         "0110010100" when "0011010", -- t[26] = 404
         "0110001110" when "0011011", -- t[27] = 398
         "0110001000" when "0011100", -- t[28] = 392
         "0110000011" when "0011101", -- t[29] = 387
         "0101111110" when "0011110", -- t[30] = 382
         "0101111001" when "0011111", -- t[31] = 377
         "0101110011" when "0100000", -- t[32] = 371
         "0101101111" when "0100001", -- t[33] = 367
         "0101101010" when "0100010", -- t[34] = 362
         "0101100101" when "0100011", -- t[35] = 357
         "0101100000" when "0100100", -- t[36] = 352
         "0101011100" when "0100101", -- t[37] = 348
         "0101010111" when "0100110", -- t[38] = 343
         "0101010011" when "0100111", -- t[39] = 339
         "0101001111" when "0101000", -- t[40] = 335
         "0101001011" when "0101001", -- t[41] = 331
         "0101000111" when "0101010", -- t[42] = 327
         "0101000011" when "0101011", -- t[43] = 323
         "0100111111" when "0101100", -- t[44] = 319
         "0100111011" when "0101101", -- t[45] = 315
         "0100110111" when "0101110", -- t[46] = 311
         "0100110011" when "0101111", -- t[47] = 307
         "0100110000" when "0110000", -- t[48] = 304
         "0100101100" when "0110001", -- t[49] = 300
         "0100101001" when "0110010", -- t[50] = 297
         "0100100101" when "0110011", -- t[51] = 293
         "0100100010" when "0110100", -- t[52] = 290
         "0100011111" when "0110101", -- t[53] = 287
         "0100011100" when "0110110", -- t[54] = 284
         "0100011001" when "0110111", -- t[55] = 281
         "0100010101" when "0111000", -- t[56] = 277
         "0100010010" when "0111001", -- t[57] = 274
         "0100001111" when "0111010", -- t[58] = 271
         "0100001101" when "0111011", -- t[59] = 269
         "0100001010" when "0111100", -- t[60] = 266
         "0100000111" when "0111101", -- t[61] = 263
         "0100000100" when "0111110", -- t[62] = 260
         "0100000001" when "0111111", -- t[63] = 257
         "0011111111" when "1000000", -- t[64] = 255
         "0011111100" when "1000001", -- t[65] = 252
         "0011111001" when "1000010", -- t[66] = 249
         "0011110111" when "1000011", -- t[67] = 247
         "0011110100" when "1000100", -- t[68] = 244
         "0011110010" when "1000101", -- t[69] = 242
         "0011110000" when "1000110", -- t[70] = 240
         "0011101101" when "1000111", -- t[71] = 237
         "0011101011" when "1001000", -- t[72] = 235
         "0011101001" when "1001001", -- t[73] = 233
         "0011100110" when "1001010", -- t[74] = 230
         "0011100100" when "1001011", -- t[75] = 228
         "0011100010" when "1001100", -- t[76] = 226
         "0011100000" when "1001101", -- t[77] = 224
         "0011011110" when "1001110", -- t[78] = 222
         "0011011100" when "1001111", -- t[79] = 220
         "0011011010" when "1010000", -- t[80] = 218
         "0011011000" when "1010001", -- t[81] = 216
         "0011010110" when "1010010", -- t[82] = 214
         "0011010100" when "1010011", -- t[83] = 212
         "0011010010" when "1010100", -- t[84] = 210
         "0011010000" when "1010101", -- t[85] = 208
         "0011001110" when "1010110", -- t[86] = 206
         "0011001100" when "1010111", -- t[87] = 204
         "0011001010" when "1011000", -- t[88] = 202
         "0011001001" when "1011001", -- t[89] = 201
         "0011000111" when "1011010", -- t[90] = 199
         "0011000101" when "1011011", -- t[91] = 197
         "0011000011" when "1011100", -- t[92] = 195
         "0011000010" when "1011101", -- t[93] = 194
         "0011000000" when "1011110", -- t[94] = 192
         "0010111110" when "1011111", -- t[95] = 190
         "0010111101" when "1100000", -- t[96] = 189
         "0010111011" when "1100001", -- t[97] = 187
         "0010111010" when "1100010", -- t[98] = 186
         "0010111000" when "1100011", -- t[99] = 184
         "0010110111" when "1100100", -- t[100] = 183
         "0010110101" when "1100101", -- t[101] = 181
         "0010110100" when "1100110", -- t[102] = 180
         "0010110010" when "1100111", -- t[103] = 178
         "0010110001" when "1101000", -- t[104] = 177
         "0010101111" when "1101001", -- t[105] = 175
         "0010101110" when "1101010", -- t[106] = 174
         "0010101100" when "1101011", -- t[107] = 172
         "0010101011" when "1101100", -- t[108] = 171
         "0010101010" when "1101101", -- t[109] = 170
         "0010101000" when "1101110", -- t[110] = 168
         "0010100111" when "1101111", -- t[111] = 167
         "0010100110" when "1110000", -- t[112] = 166
         "0010100101" when "1110001", -- t[113] = 165
         "0010100011" when "1110010", -- t[114] = 163
         "0010100010" when "1110011", -- t[115] = 162
         "0010100001" when "1110100", -- t[116] = 161
         "0010100000" when "1110101", -- t[117] = 160
         "0010011110" when "1110110", -- t[118] = 158
         "0010011101" when "1110111", -- t[119] = 157
         "0010011100" when "1111000", -- t[120] = 156
         "0010011011" when "1111001", -- t[121] = 155
         "0010011010" when "1111010", -- t[122] = 154
         "0010011001" when "1111011", -- t[123] = 153
         "0010011000" when "1111100", -- t[124] = 152
         "0010010110" when "1111101", -- t[125] = 150
         "0010010101" when "1111110", -- t[126] = 149
         "0010010100" when "1111111", -- t[127] = 148
         "----------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 7; beta_1 = 7; lambda_1 = 7;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 7; rho_1,1 = 0; sigma_1,1 = 7; wO_1,1 = 10.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_14_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of fp_log_log_14_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(5 downto 0);
  signal s      : std_logic_vector(6 downto 0);
  component fp_log_log_14_t1_pow is
    port ( x : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(5 downto 0);
  signal k_1    : std_logic_vector(9 downto 0);
  signal r0_1   : std_logic_vector(17 downto 0);
  signal r_1    : std_logic_vector(16 downto 0);
  component fp_log_log_14_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;
begin
  sign <= not b(6);
  b0 <= b(5 downto 0) xor (5 downto 0 => sign);

  pow : fp_log_log_14_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(6);
  s_1 <= s(5 downto 0) xor (5 downto 0 => sign_1);
  t_1 : fp_log_log_14_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(9 downto 0) <=
    r0_1(17 downto 8) xor (17 downto 8 => (not (sign xor sign_1)));
  r_1(16 downto 10) <= (16 downto 10 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_14 is
  port ( x : in  std_logic_vector(13 downto 0);
         r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of fp_log_log_14 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(16 downto 0);
  component fp_log_log_14_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(16 downto 0) );
  end component;

  signal a_1 : std_logic_vector(6 downto 0);
  signal b_1 : std_logic_vector(6 downto 0);
  signal r_1 : std_logic_vector(16 downto 0);
  component fp_log_log_14_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(16 downto 0) );
  end component;

begin
  a_0 <= x(13 downto 7);
  t_0 : fp_log_log_14_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(13 downto 7);
  b_1 <= x(6 downto 0);
  t_1 : fp_log_log_14_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  r <= r_0 + r_1;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 15; wO = 15.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 8;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 7; beta_1 = 8;
--   T_2 (ROM):     alpha_2 = 2; beta_2 = 2.
-- Guard bits: g = 4.
-- Command line: logfp 15 15 2   rom 7 0   pm 7 8  ah 8 8 8  1 1  7 6 0  4 2 6   rom 2 2


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 20.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_15_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_15_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(19 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110000110101101001" when "0000000", -- t[0] = 724329
          "10101111101000100111" when "0000001", -- t[1] = 719399
          "10101110011101000010" when "0000010", -- t[2] = 714562
          "10101101010010111000" when "0000011", -- t[3] = 709816
          "10101100001010000110" when "0000100", -- t[4] = 705158
          "10101011000010101010" when "0000101", -- t[5] = 700586
          "10101001111100100000" when "0000110", -- t[6] = 696096
          "10101000110111100111" when "0000111", -- t[7] = 691687
          "10100111110011111011" when "0001000", -- t[8] = 687355
          "10100110110001011010" when "0001001", -- t[9] = 683098
          "10100101110000000011" when "0001010", -- t[10] = 678915
          "10100100101111110010" when "0001011", -- t[11] = 674802
          "10100011110000100110" when "0001100", -- t[12] = 670758
          "10100010110010011110" when "0001101", -- t[13] = 666782
          "10100001110101010110" when "0001110", -- t[14] = 662870
          "10100000111001001110" when "0001111", -- t[15] = 659022
          "10011111111110000011" when "0010000", -- t[16] = 655235
          "10011111000011110100" when "0010001", -- t[17] = 651508
          "10011110001010100000" when "0010010", -- t[18] = 647840
          "10011101010010000100" when "0010011", -- t[19] = 644228
          "10011100011010011111" when "0010100", -- t[20] = 640671
          "10011011100011110000" when "0010101", -- t[21] = 637168
          "10011010101101110110" when "0010110", -- t[22] = 633718
          "10011001111000101111" when "0010111", -- t[23] = 630319
          "10011001000100011001" when "0011000", -- t[24] = 626969
          "10011000010000110100" when "0011001", -- t[25] = 623668
          "10010111011101111111" when "0011010", -- t[26] = 620415
          "10010110101011111000" when "0011011", -- t[27] = 617208
          "10010101111010011110" when "0011100", -- t[28] = 614046
          "10010101001001110000" when "0011101", -- t[29] = 610928
          "10010100011001101100" when "0011110", -- t[30] = 607852
          "10010011101010010011" when "0011111", -- t[31] = 604819
          "10010010111011100110" when "0100000", -- t[32] = 601830
          "10010010001101011110" when "0100001", -- t[33] = 598878
          "10010001011111111110" when "0100010", -- t[34] = 595966
          "10010000110011000011" when "0100011", -- t[35] = 593091
          "10010000000110101110" when "0100100", -- t[36] = 590254
          "10001111011010111110" when "0100101", -- t[37] = 587454
          "10001110101111110010" when "0100110", -- t[38] = 584690
          "10001110000101001000" when "0100111", -- t[39] = 581960
          "10001101011011000010" when "0101000", -- t[40] = 579266
          "10001100110001011100" when "0101001", -- t[41] = 576604
          "10001100001000011000" when "0101010", -- t[42] = 573976
          "10001011011111110011" when "0101011", -- t[43] = 571379
          "10001010110111101111" when "0101100", -- t[44] = 568815
          "10001010010000001001" when "0101101", -- t[45] = 566281
          "10001001101001000001" when "0101110", -- t[46] = 563777
          "10001001000010010111" when "0101111", -- t[47] = 561303
          "10001000011100001011" when "0110000", -- t[48] = 558859
          "10000111110110011010" when "0110001", -- t[49] = 556442
          "10000111010001000110" when "0110010", -- t[50] = 554054
          "10000110101100001101" when "0110011", -- t[51] = 551693
          "10000110000111101111" when "0110100", -- t[52] = 549359
          "10000101100011101011" when "0110101", -- t[53] = 547051
          "10000101000000000001" when "0110110", -- t[54] = 544769
          "10000100011100110001" when "0110111", -- t[55] = 542513
          "10000011111001111001" when "0111000", -- t[56] = 540281
          "10000011010111011010" when "0111001", -- t[57] = 538074
          "10000010110101010011" when "0111010", -- t[58] = 535891
          "10000010010011100011" when "0111011", -- t[59] = 533731
          "10000001110010001010" when "0111100", -- t[60] = 531594
          "10000001010001001001" when "0111101", -- t[61] = 529481
          "10000000110000011101" when "0111110", -- t[62] = 527389
          "10000000010000000111" when "0111111", -- t[63] = 525319
          "01111111110000001000" when "1000000", -- t[64] = 523272
          "01111111010000011110" when "1000001", -- t[65] = 521246
          "01111110110001000111" when "1000010", -- t[66] = 519239
          "01111110010010000110" when "1000011", -- t[67] = 517254
          "01111101110011011000" when "1000100", -- t[68] = 515288
          "01111101010100111110" when "1000101", -- t[69] = 513342
          "01111100110110111000" when "1000110", -- t[70] = 511416
          "01111100011001000100" when "1000111", -- t[71] = 509508
          "01111011111011100011" when "1001000", -- t[72] = 507619
          "01111011011110010101" when "1001001", -- t[73] = 505749
          "01111011000001011001" when "1001010", -- t[74] = 503897
          "01111010100100101111" when "1001011", -- t[75] = 502063
          "01111010001000010110" when "1001100", -- t[76] = 500246
          "01111001101100001111" when "1001101", -- t[77] = 498447
          "01111001010000011001" when "1001110", -- t[78] = 496665
          "01111000110100110011" when "1001111", -- t[79] = 494899
          "01111000011001011110" when "1010000", -- t[80] = 493150
          "01110111111110011001" when "1010001", -- t[81] = 491417
          "01110111100011100101" when "1010010", -- t[82] = 489701
          "01110111001000111111" when "1010011", -- t[83] = 487999
          "01110110101110101010" when "1010100", -- t[84] = 486314
          "01110110010100100011" when "1010101", -- t[85] = 484643
          "01110101111010101100" when "1010110", -- t[86] = 482988
          "01110101100001000011" when "1010111", -- t[87] = 481347
          "01110101000111101001" when "1011000", -- t[88] = 479721
          "01110100101110011110" when "1011001", -- t[89] = 478110
          "01110100010101100000" when "1011010", -- t[90] = 476512
          "01110011111100110001" when "1011011", -- t[91] = 474929
          "01110011100100001111" when "1011100", -- t[92] = 473359
          "01110011001011111011" when "1011101", -- t[93] = 471803
          "01110010110011110100" when "1011110", -- t[94] = 470260
          "01110010011011111010" when "1011111", -- t[95] = 468730
          "01110010000100001110" when "1100000", -- t[96] = 467214
          "01110001101100101110" when "1100001", -- t[97] = 465710
          "01110001010101011010" when "1100010", -- t[98] = 464218
          "01110000111110010011" when "1100011", -- t[99] = 462739
          "01110000100111011001" when "1100100", -- t[100] = 461273
          "01110000010000101010" when "1100101", -- t[101] = 459818
          "01101111111010000111" when "1100110", -- t[102] = 458375
          "01101111100011110001" when "1100111", -- t[103] = 456945
          "01101111001101100101" when "1101000", -- t[104] = 455525
          "01101110110111100101" when "1101001", -- t[105] = 454117
          "01101110100001110001" when "1101010", -- t[106] = 452721
          "01101110001100000111" when "1101011", -- t[107] = 451335
          "01101101110110101001" when "1101100", -- t[108] = 449961
          "01101101100001010101" when "1101101", -- t[109] = 448597
          "01101101001100001100" when "1101110", -- t[110] = 447244
          "01101100110111001110" when "1101111", -- t[111] = 445902
          "01101100100010011010" when "1110000", -- t[112] = 444570
          "01101100001101110000" when "1110001", -- t[113] = 443248
          "01101011111001010001" when "1110010", -- t[114] = 441937
          "01101011100100111011" when "1110011", -- t[115] = 440635
          "01101011010000110000" when "1110100", -- t[116] = 439344
          "01101010111100101110" when "1110101", -- t[117] = 438062
          "01101010101000110110" when "1110110", -- t[118] = 436790
          "01101010010101001000" when "1110111", -- t[119] = 435528
          "01101010000001100010" when "1111000", -- t[120] = 434274
          "01101001101110000111" when "1111001", -- t[121] = 433031
          "01101001011010110100" when "1111010", -- t[122] = 431796
          "01101001000111101010" when "1111011", -- t[123] = 430570
          "01101000110100101010" when "1111100", -- t[124] = 429354
          "01101000100001110010" when "1111101", -- t[125] = 428146
          "01101000001111000011" when "1111110", -- t[126] = 426947
          "01100111111100011101" when "1111111", -- t[127] = 425757
          "--------------------" when others;

  r(19 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 8; mu_1 = 8; lambda_1 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_15_t1_pow is
  port ( x : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_log_log_15_t1_pow is
  signal pp0 : std_logic_vector(6 downto 0);
  signal r0 : std_logic_vector(6 downto 0);
begin
  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(6 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 7; wO_1,1 = 13.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_15_t1_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of fp_log_log_15_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "1001101110011" when "0000000", -- t[0] = 4979
         "1001100010011" when "0000001", -- t[1] = 4883
         "1001010110111" when "0000010", -- t[2] = 4791
         "1001001011101" when "0000011", -- t[3] = 4701
         "1001000000110" when "0000100", -- t[4] = 4614
         "1000110110011" when "0000101", -- t[5] = 4531
         "1000101100001" when "0000110", -- t[6] = 4449
         "1000100010010" when "0000111", -- t[7] = 4370
         "1000011000110" when "0001000", -- t[8] = 4294
         "1000001111100" when "0001001", -- t[9] = 4220
         "1000000110100" when "0001010", -- t[10] = 4148
         "0111111101110" when "0001011", -- t[11] = 4078
         "0111110101010" when "0001100", -- t[12] = 4010
         "0111101101000" when "0001101", -- t[13] = 3944
         "0111100101000" when "0001110", -- t[14] = 3880
         "0111011101001" when "0001111", -- t[15] = 3817
         "0111010101100" when "0010000", -- t[16] = 3756
         "0111001110001" when "0010001", -- t[17] = 3697
         "0111000111000" when "0010010", -- t[18] = 3640
         "0111000000000" when "0010011", -- t[19] = 3584
         "0110111001001" when "0010100", -- t[20] = 3529
         "0110110010100" when "0010101", -- t[21] = 3476
         "0110101100001" when "0010110", -- t[22] = 3425
         "0110100101110" when "0010111", -- t[23] = 3374
         "0110011111101" when "0011000", -- t[24] = 3325
         "0110011001101" when "0011001", -- t[25] = 3277
         "0110010011110" when "0011010", -- t[26] = 3230
         "0110001110000" when "0011011", -- t[27] = 3184
         "0110001000100" when "0011100", -- t[28] = 3140
         "0110000011000" when "0011101", -- t[29] = 3096
         "0101111101110" when "0011110", -- t[30] = 3054
         "0101111000100" when "0011111", -- t[31] = 3012
         "0101110011100" when "0100000", -- t[32] = 2972
         "0101101110100" when "0100001", -- t[33] = 2932
         "0101101001101" when "0100010", -- t[34] = 2893
         "0101100100111" when "0100011", -- t[35] = 2855
         "0101100000010" when "0100100", -- t[36] = 2818
         "0101011011110" when "0100101", -- t[37] = 2782
         "0101010111011" when "0100110", -- t[38] = 2747
         "0101010011000" when "0100111", -- t[39] = 2712
         "0101001110110" when "0101000", -- t[40] = 2678
         "0101001010101" when "0101001", -- t[41] = 2645
         "0101000110100" when "0101010", -- t[42] = 2612
         "0101000010100" when "0101011", -- t[43] = 2580
         "0100111110101" when "0101100", -- t[44] = 2549
         "0100111010111" when "0101101", -- t[45] = 2519
         "0100110111001" when "0101110", -- t[46] = 2489
         "0100110011011" when "0101111", -- t[47] = 2459
         "0100101111110" when "0110000", -- t[48] = 2430
         "0100101100010" when "0110001", -- t[49] = 2402
         "0100101000111" when "0110010", -- t[50] = 2375
         "0100100101011" when "0110011", -- t[51] = 2347
         "0100100010001" when "0110100", -- t[52] = 2321
         "0100011110111" when "0110101", -- t[53] = 2295
         "0100011011101" when "0110110", -- t[54] = 2269
         "0100011000100" when "0110111", -- t[55] = 2244
         "0100010101011" when "0111000", -- t[56] = 2219
         "0100010010011" when "0111001", -- t[57] = 2195
         "0100001111011" when "0111010", -- t[58] = 2171
         "0100001100100" when "0111011", -- t[59] = 2148
         "0100001001101" when "0111100", -- t[60] = 2125
         "0100000110111" when "0111101", -- t[61] = 2103
         "0100000100000" when "0111110", -- t[62] = 2080
         "0100000001011" when "0111111", -- t[63] = 2059
         "0011111110101" when "1000000", -- t[64] = 2037
         "0011111100000" when "1000001", -- t[65] = 2016
         "0011111001100" when "1000010", -- t[66] = 1996
         "0011110111000" when "1000011", -- t[67] = 1976
         "0011110100100" when "1000100", -- t[68] = 1956
         "0011110010000" when "1000101", -- t[69] = 1936
         "0011101111101" when "1000110", -- t[70] = 1917
         "0011101101010" when "1000111", -- t[71] = 1898
         "0011101010111" when "1001000", -- t[72] = 1879
         "0011101000101" when "1001001", -- t[73] = 1861
         "0011100110011" when "1001010", -- t[74] = 1843
         "0011100100001" when "1001011", -- t[75] = 1825
         "0011100010000" when "1001100", -- t[76] = 1808
         "0011011111111" when "1001101", -- t[77] = 1791
         "0011011101110" when "1001110", -- t[78] = 1774
         "0011011011101" when "1001111", -- t[79] = 1757
         "0011011001101" when "1010000", -- t[80] = 1741
         "0011010111101" when "1010001", -- t[81] = 1725
         "0011010101101" when "1010010", -- t[82] = 1709
         "0011010011101" when "1010011", -- t[83] = 1693
         "0011010001110" when "1010100", -- t[84] = 1678
         "0011001111111" when "1010101", -- t[85] = 1663
         "0011001110000" when "1010110", -- t[86] = 1648
         "0011001100001" when "1010111", -- t[87] = 1633
         "0011001010011" when "1011000", -- t[88] = 1619
         "0011001000101" when "1011001", -- t[89] = 1605
         "0011000110110" when "1011010", -- t[90] = 1590
         "0011000101001" when "1011011", -- t[91] = 1577
         "0011000011011" when "1011100", -- t[92] = 1563
         "0011000001110" when "1011101", -- t[93] = 1550
         "0011000000000" when "1011110", -- t[94] = 1536
         "0010111110011" when "1011111", -- t[95] = 1523
         "0010111100110" when "1100000", -- t[96] = 1510
         "0010111011010" when "1100001", -- t[97] = 1498
         "0010111001101" when "1100010", -- t[98] = 1485
         "0010111000001" when "1100011", -- t[99] = 1473
         "0010110110101" when "1100100", -- t[100] = 1461
         "0010110101001" when "1100101", -- t[101] = 1449
         "0010110011101" when "1100110", -- t[102] = 1437
         "0010110010001" when "1100111", -- t[103] = 1425
         "0010110000110" when "1101000", -- t[104] = 1414
         "0010101111010" when "1101001", -- t[105] = 1402
         "0010101101111" when "1101010", -- t[106] = 1391
         "0010101100100" when "1101011", -- t[107] = 1380
         "0010101011001" when "1101100", -- t[108] = 1369
         "0010101001110" when "1101101", -- t[109] = 1358
         "0010101000100" when "1101110", -- t[110] = 1348
         "0010100111001" when "1101111", -- t[111] = 1337
         "0010100101111" when "1110000", -- t[112] = 1327
         "0010100100101" when "1110001", -- t[113] = 1317
         "0010100011010" when "1110010", -- t[114] = 1306
         "0010100010000" when "1110011", -- t[115] = 1296
         "0010100000111" when "1110100", -- t[116] = 1287
         "0010011111101" when "1110101", -- t[117] = 1277
         "0010011110011" when "1110110", -- t[118] = 1267
         "0010011101010" when "1110111", -- t[119] = 1258
         "0010011100000" when "1111000", -- t[120] = 1248
         "0010011010111" when "1111001", -- t[121] = 1239
         "0010011001110" when "1111010", -- t[122] = 1230
         "0010011000101" when "1111011", -- t[123] = 1221
         "0010010111100" when "1111100", -- t[124] = 1212
         "0010010110011" when "1111101", -- t[125] = 1203
         "0010010101011" when "1111110", -- t[126] = 1195
         "0010010100010" when "1111111", -- t[127] = 1186
         "-------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_2.
-- Decomposition:
--   alpha_1,2 = 4; sigma'_1,2 = 1; wO_1,2 = 5.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_15_t1_t2 is
  port ( a : in  std_logic_vector(3 downto 0);
         s : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of fp_log_log_15_t1_t2 is
  signal x : std_logic_vector(4 downto 0);
begin
  x <= a & s;

  with x select
    r <= "01001" when "00000", -- t[0] = 9
         "11011" when "00001", -- t[1] = 27
         "00111" when "00010", -- t[2] = 7
         "10111" when "00011", -- t[3] = 23
         "00110" when "00100", -- t[4] = 6
         "10100" when "00101", -- t[5] = 20
         "00110" when "00110", -- t[6] = 6
         "10010" when "00111", -- t[7] = 18
         "00101" when "01000", -- t[8] = 5
         "10000" when "01001", -- t[9] = 16
         "00101" when "01010", -- t[10] = 5
         "01111" when "01011", -- t[11] = 15
         "00100" when "01100", -- t[12] = 4
         "01101" when "01101", -- t[13] = 13
         "00100" when "01110", -- t[14] = 4
         "01100" when "01111", -- t[15] = 12
         "00011" when "10000", -- t[16] = 3
         "01011" when "10001", -- t[17] = 11
         "00011" when "10010", -- t[18] = 3
         "01010" when "10011", -- t[19] = 10
         "00011" when "10100", -- t[20] = 3
         "01001" when "10101", -- t[21] = 9
         "00011" when "10110", -- t[22] = 3
         "01001" when "10111", -- t[23] = 9
         "00010" when "11000", -- t[24] = 2
         "01000" when "11001", -- t[25] = 8
         "00010" when "11010", -- t[26] = 2
         "01000" when "11011", -- t[27] = 8
         "00010" when "11100", -- t[28] = 2
         "00111" when "11101", -- t[29] = 7
         "00010" when "11110", -- t[30] = 2
         "00111" when "11111", -- t[31] = 7
         "-----" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 7; beta_1 = 8; lambda_1 = 8;  m_1 = 2;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 7; rho_1,1 = 0; sigma_1,1 = 6; wO_1,1 = 13;
--   Q_1,2 (ROM):  alpha_1,2 = 4; rho_1,2 = 6; sigma_1,2 = 2; wO_1,2 = 5.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_15_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_15_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(6 downto 0);
  signal s      : std_logic_vector(7 downto 0);
  component fp_log_log_15_t1_pow is
    port ( x : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(4 downto 0);
  signal k_1    : std_logic_vector(12 downto 0);
  signal r0_1   : std_logic_vector(19 downto 0);
  signal r_1    : std_logic_vector(19 downto 0);
  component fp_log_log_15_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  signal a_2    : std_logic_vector(3 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(0 downto 0);
  signal r0_2   : std_logic_vector(4 downto 0);
  signal r_2    : std_logic_vector(19 downto 0);
  component fp_log_log_15_t1_t2 is
    port ( a : in  std_logic_vector(3 downto 0);
           s : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;
begin
  sign <= not b(7);
  b0 <= b(6 downto 0) xor (6 downto 0 => sign);

  pow : fp_log_log_15_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(7);
  s_1 <= s(6 downto 2) xor (6 downto 2 => sign_1);
  t_1 : fp_log_log_15_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(12 downto 0) <=
    r0_1(19 downto 7) xor (19 downto 7 => (not (sign xor sign_1)));
  r_1(19 downto 13) <= (19 downto 13 => (not (sign xor sign_1)));

  a_2 <= a(6 downto 3);
  sign_2 <= not s(1);
  s_2 <= s(0 downto 0) xor (0 downto 0 => sign_2);
  t_2 : fp_log_log_15_t1_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(4 downto 0) <=
    r0_2 xor (4 downto 0 => (not (sign xor sign_2)));
  r_2(19 downto 5) <= (19 downto 5 => (not (sign xor sign_2)));

  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- TermROM instance for order-2 term.
-- Decomposition:
--   alpha_2 = 2; beta_2 = 2 (1+1); wO_2 = 3.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_15_t2 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_15_t2 is
  signal sign : std_logic;
  signal b0   : std_logic_vector(0 downto 0);
  signal x0   : std_logic_vector(2 downto 0);
  signal r0   : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  b0 <= b(0 downto 0) xor (0 downto 0 => sign);
  x0 <= a & b0;

  with x0 select
    r0 <= "001" when "000", -- t[0] = 1
          "101" when "001", -- t[1] = 5
          "000" when "010", -- t[2] = 0
          "010" when "011", -- t[3] = 2
          "000" when "100", -- t[4] = 0
          "001" when "101", -- t[5] = 1
          "000" when "110", -- t[6] = 0
          "000" when "111", -- t[7] = 0
          "---" when others;

  r(2 downto 0) <= r0;
  r(19 downto 3) <= (19 downto 3 => ('0'));
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_15 is
  port ( x : in  std_logic_vector(14 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_15 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(19 downto 0);
  component fp_log_log_15_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

  signal a_1 : std_logic_vector(6 downto 0);
  signal b_1 : std_logic_vector(7 downto 0);
  signal r_1 : std_logic_vector(19 downto 0);
  component fp_log_log_15_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

  signal a_2 : std_logic_vector(1 downto 0);
  signal b_2 : std_logic_vector(1 downto 0);
  signal r_2 : std_logic_vector(19 downto 0);
  component fp_log_log_15_t2 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

begin
  a_0 <= x(14 downto 8);
  t_0 : fp_log_log_15_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(14 downto 8);
  b_1 <= x(7 downto 0);
  t_1 : fp_log_log_15_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(14 downto 13);
  b_2 <= x(7 downto 6);
  t_2 : fp_log_log_15_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 16; wO = 16.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 9;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 7; beta_1 = 9;
--   T_2 (ROM):     alpha_2 = 3; beta_2 = 4.
-- Guard bits: g = 3.
-- Command line: logfp 16 16 2   rom 7 0   pm 7 9  ah 9 9 9  1 0  7 9 0   rom 3 4


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 20.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_16_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_16_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(19 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110000110101100011" when "0000000", -- t[0] = 724323
          "10101111101000100001" when "0000001", -- t[1] = 719393
          "10101110011100111100" when "0000010", -- t[2] = 714556
          "10101101010010110010" when "0000011", -- t[3] = 709810
          "10101100001010000001" when "0000100", -- t[4] = 705153
          "10101011000010100100" when "0000101", -- t[5] = 700580
          "10101001111100011011" when "0000110", -- t[6] = 696091
          "10101000110111100001" when "0000111", -- t[7] = 691681
          "10100111110011110101" when "0001000", -- t[8] = 687349
          "10100110110001010100" when "0001001", -- t[9] = 683092
          "10100101101111111101" when "0001010", -- t[10] = 678909
          "10100100101111101101" when "0001011", -- t[11] = 674797
          "10100011110000100001" when "0001100", -- t[12] = 670753
          "10100010110010011001" when "0001101", -- t[13] = 666777
          "10100001110101010001" when "0001110", -- t[14] = 662865
          "10100000111001001001" when "0001111", -- t[15] = 659017
          "10011111111110000001" when "0010000", -- t[16] = 655233
          "10011111000011110010" when "0010001", -- t[17] = 651506
          "10011110001010011101" when "0010010", -- t[18] = 647837
          "10011101010010000001" when "0010011", -- t[19] = 644225
          "10011100011010011101" when "0010100", -- t[20] = 640669
          "10011011100011101110" when "0010101", -- t[21] = 637166
          "10011010101101110100" when "0010110", -- t[22] = 633716
          "10011001111000101100" when "0010111", -- t[23] = 630316
          "10011001000100010111" when "0011000", -- t[24] = 626967
          "10011000010000110010" when "0011001", -- t[25] = 623666
          "10010111011101111100" when "0011010", -- t[26] = 620412
          "10010110101011110101" when "0011011", -- t[27] = 617205
          "10010101111010011011" when "0011100", -- t[28] = 614043
          "10010101001001101101" when "0011101", -- t[29] = 610925
          "10010100011001101010" when "0011110", -- t[30] = 607850
          "10010011101010010001" when "0011111", -- t[31] = 604817
          "10010010111011100011" when "0100000", -- t[32] = 601827
          "10010010001101011011" when "0100001", -- t[33] = 598875
          "10010001011111111010" when "0100010", -- t[34] = 595962
          "10010000110011000000" when "0100011", -- t[35] = 593088
          "10010000000110101011" when "0100100", -- t[36] = 590251
          "10001111011010111011" when "0100101", -- t[37] = 587451
          "10001110101111101110" when "0100110", -- t[38] = 584686
          "10001110000101000101" when "0100111", -- t[39] = 581957
          "10001101011010111110" when "0101000", -- t[40] = 579262
          "10001100110001011001" when "0101001", -- t[41] = 576601
          "10001100001000010100" when "0101010", -- t[42] = 573972
          "10001011011111110000" when "0101011", -- t[43] = 571376
          "10001010110111101011" when "0101100", -- t[44] = 568811
          "10001010010000000101" when "0101101", -- t[45] = 566277
          "10001001101000111110" when "0101110", -- t[46] = 563774
          "10001001000010010100" when "0101111", -- t[47] = 561300
          "10001000011100001000" when "0110000", -- t[48] = 558856
          "10000111110110011000" when "0110001", -- t[49] = 556440
          "10000111010001000100" when "0110010", -- t[50] = 554052
          "10000110101100001011" when "0110011", -- t[51] = 551691
          "10000110000111101101" when "0110100", -- t[52] = 549357
          "10000101100011101001" when "0110101", -- t[53] = 547049
          "10000100111111111111" when "0110110", -- t[54] = 544767
          "10000100011100101110" when "0110111", -- t[55] = 542510
          "10000011111001110111" when "0111000", -- t[56] = 540279
          "10000011010111011000" when "0111001", -- t[57] = 538072
          "10000010110101010000" when "0111010", -- t[58] = 535888
          "10000010010011100001" when "0111011", -- t[59] = 533729
          "10000001110010001000" when "0111100", -- t[60] = 531592
          "10000001010001000110" when "0111101", -- t[61] = 529478
          "10000000110000011011" when "0111110", -- t[62] = 527387
          "10000000010000000101" when "0111111", -- t[63] = 525317
          "01111111110000000110" when "1000000", -- t[64] = 523270
          "01111111010000011011" when "1000001", -- t[65] = 521243
          "01111110110001000101" when "1000010", -- t[66] = 519237
          "01111110010010000011" when "1000011", -- t[67] = 517251
          "01111101110011010101" when "1000100", -- t[68] = 515285
          "01111101010100111100" when "1000101", -- t[69] = 513340
          "01111100110110110101" when "1000110", -- t[70] = 511413
          "01111100011001000010" when "1000111", -- t[71] = 509506
          "01111011111011100001" when "1001000", -- t[72] = 507617
          "01111011011110010011" when "1001001", -- t[73] = 505747
          "01111011000001010111" when "1001010", -- t[74] = 503895
          "01111010100100101101" when "1001011", -- t[75] = 502061
          "01111010001000010100" when "1001100", -- t[76] = 500244
          "01111001101100001101" when "1001101", -- t[77] = 498445
          "01111001010000010110" when "1001110", -- t[78] = 496662
          "01111000110100110001" when "1001111", -- t[79] = 494897
          "01111000011001011100" when "1010000", -- t[80] = 493148
          "01110111111110010111" when "1010001", -- t[81] = 491415
          "01110111100011100011" when "1010010", -- t[82] = 489699
          "01110111001000111101" when "1010011", -- t[83] = 487997
          "01110110101110101000" when "1010100", -- t[84] = 486312
          "01110110010100100001" when "1010101", -- t[85] = 484641
          "01110101111010101010" when "1010110", -- t[86] = 482986
          "01110101100001000010" when "1010111", -- t[87] = 481346
          "01110101000111101000" when "1011000", -- t[88] = 479720
          "01110100101110011100" when "1011001", -- t[89] = 478108
          "01110100010101011110" when "1011010", -- t[90] = 476510
          "01110011111100101111" when "1011011", -- t[91] = 474927
          "01110011100100001101" when "1011100", -- t[92] = 473357
          "01110011001011111001" when "1011101", -- t[93] = 471801
          "01110010110011110010" when "1011110", -- t[94] = 470258
          "01110010011011111000" when "1011111", -- t[95] = 468728
          "01110010000100001100" when "1100000", -- t[96] = 467212
          "01110001101100101100" when "1100001", -- t[97] = 465708
          "01110001010101011000" when "1100010", -- t[98] = 464216
          "01110000111110010001" when "1100011", -- t[99] = 462737
          "01110000100111010111" when "1100100", -- t[100] = 461271
          "01110000010000101000" when "1100101", -- t[101] = 459816
          "01101111111010000101" when "1100110", -- t[102] = 458373
          "01101111100011101111" when "1100111", -- t[103] = 456943
          "01101111001101100011" when "1101000", -- t[104] = 455523
          "01101110110111100011" when "1101001", -- t[105] = 454115
          "01101110100001101111" when "1101010", -- t[106] = 452719
          "01101110001100000101" when "1101011", -- t[107] = 451333
          "01101101110110100111" when "1101100", -- t[108] = 449959
          "01101101100001010011" when "1101101", -- t[109] = 448595
          "01101101001100001010" when "1101110", -- t[110] = 447242
          "01101100110111001100" when "1101111", -- t[111] = 445900
          "01101100100010011000" when "1110000", -- t[112] = 444568
          "01101100001101101111" when "1110001", -- t[113] = 443247
          "01101011111001001111" when "1110010", -- t[114] = 441935
          "01101011100100111010" when "1110011", -- t[115] = 440634
          "01101011010000101110" when "1110100", -- t[116] = 439342
          "01101010111100101101" when "1110101", -- t[117] = 438061
          "01101010101000110100" when "1110110", -- t[118] = 436788
          "01101010010101000110" when "1110111", -- t[119] = 435526
          "01101010000001100001" when "1111000", -- t[120] = 434273
          "01101001101110000101" when "1111001", -- t[121] = 433029
          "01101001011010110010" when "1111010", -- t[122] = 431794
          "01101001000111101001" when "1111011", -- t[123] = 430569
          "01101000110100101000" when "1111100", -- t[124] = 429352
          "01101000100001110000" when "1111101", -- t[125] = 428144
          "01101000001111000001" when "1111110", -- t[126] = 426945
          "01100111111100011011" when "1111111", -- t[127] = 425755
          "--------------------" when others;

  r(19 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 9; mu_1 = 9; lambda_1 = 9.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_16_t1_pow is
  port ( x : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of fp_log_log_16_t1_pow is
  signal pp0 : std_logic_vector(7 downto 0);
  signal r0 : std_logic_vector(7 downto 0);
begin
  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(7 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 7; wO_1,1 = 13.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_16_t1_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of fp_log_log_16_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "1001101110011" when "0000000", -- t[0] = 4979
         "1001100010011" when "0000001", -- t[1] = 4883
         "1001010110111" when "0000010", -- t[2] = 4791
         "1001001011101" when "0000011", -- t[3] = 4701
         "1001000000110" when "0000100", -- t[4] = 4614
         "1000110110010" when "0000101", -- t[5] = 4530
         "1000101100001" when "0000110", -- t[6] = 4449
         "1000100010010" when "0000111", -- t[7] = 4370
         "1000011000110" when "0001000", -- t[8] = 4294
         "1000001111100" when "0001001", -- t[9] = 4220
         "1000000110100" when "0001010", -- t[10] = 4148
         "0111111101110" when "0001011", -- t[11] = 4078
         "0111110101010" when "0001100", -- t[12] = 4010
         "0111101101000" when "0001101", -- t[13] = 3944
         "0111100100111" when "0001110", -- t[14] = 3879
         "0111011101001" when "0001111", -- t[15] = 3817
         "0111010101100" when "0010000", -- t[16] = 3756
         "0111001110001" when "0010001", -- t[17] = 3697
         "0111000111000" when "0010010", -- t[18] = 3640
         "0111000000000" when "0010011", -- t[19] = 3584
         "0110111001001" when "0010100", -- t[20] = 3529
         "0110110010100" when "0010101", -- t[21] = 3476
         "0110101100001" when "0010110", -- t[22] = 3425
         "0110100101110" when "0010111", -- t[23] = 3374
         "0110011111101" when "0011000", -- t[24] = 3325
         "0110011001101" when "0011001", -- t[25] = 3277
         "0110010011110" when "0011010", -- t[26] = 3230
         "0110001110000" when "0011011", -- t[27] = 3184
         "0110001000100" when "0011100", -- t[28] = 3140
         "0110000011000" when "0011101", -- t[29] = 3096
         "0101111101110" when "0011110", -- t[30] = 3054
         "0101111000100" when "0011111", -- t[31] = 3012
         "0101110011100" when "0100000", -- t[32] = 2972
         "0101101110100" when "0100001", -- t[33] = 2932
         "0101101001101" when "0100010", -- t[34] = 2893
         "0101100100111" when "0100011", -- t[35] = 2855
         "0101100000010" when "0100100", -- t[36] = 2818
         "0101011011110" when "0100101", -- t[37] = 2782
         "0101010111011" when "0100110", -- t[38] = 2747
         "0101010011000" when "0100111", -- t[39] = 2712
         "0101001110110" when "0101000", -- t[40] = 2678
         "0101001010101" when "0101001", -- t[41] = 2645
         "0101000110100" when "0101010", -- t[42] = 2612
         "0101000010100" when "0101011", -- t[43] = 2580
         "0100111110101" when "0101100", -- t[44] = 2549
         "0100111010111" when "0101101", -- t[45] = 2519
         "0100110111001" when "0101110", -- t[46] = 2489
         "0100110011011" when "0101111", -- t[47] = 2459
         "0100101111110" when "0110000", -- t[48] = 2430
         "0100101100010" when "0110001", -- t[49] = 2402
         "0100101000111" when "0110010", -- t[50] = 2375
         "0100100101011" when "0110011", -- t[51] = 2347
         "0100100010001" when "0110100", -- t[52] = 2321
         "0100011110111" when "0110101", -- t[53] = 2295
         "0100011011101" when "0110110", -- t[54] = 2269
         "0100011000100" when "0110111", -- t[55] = 2244
         "0100010101011" when "0111000", -- t[56] = 2219
         "0100010010011" when "0111001", -- t[57] = 2195
         "0100001111011" when "0111010", -- t[58] = 2171
         "0100001100100" when "0111011", -- t[59] = 2148
         "0100001001101" when "0111100", -- t[60] = 2125
         "0100000110111" when "0111101", -- t[61] = 2103
         "0100000100000" when "0111110", -- t[62] = 2080
         "0100000001011" when "0111111", -- t[63] = 2059
         "0011111110101" when "1000000", -- t[64] = 2037
         "0011111100000" when "1000001", -- t[65] = 2016
         "0011111001100" when "1000010", -- t[66] = 1996
         "0011110111000" when "1000011", -- t[67] = 1976
         "0011110100100" when "1000100", -- t[68] = 1956
         "0011110010000" when "1000101", -- t[69] = 1936
         "0011101111101" when "1000110", -- t[70] = 1917
         "0011101101010" when "1000111", -- t[71] = 1898
         "0011101010111" when "1001000", -- t[72] = 1879
         "0011101000101" when "1001001", -- t[73] = 1861
         "0011100110011" when "1001010", -- t[74] = 1843
         "0011100100001" when "1001011", -- t[75] = 1825
         "0011100010000" when "1001100", -- t[76] = 1808
         "0011011111111" when "1001101", -- t[77] = 1791
         "0011011101110" when "1001110", -- t[78] = 1774
         "0011011011101" when "1001111", -- t[79] = 1757
         "0011011001101" when "1010000", -- t[80] = 1741
         "0011010111101" when "1010001", -- t[81] = 1725
         "0011010101101" when "1010010", -- t[82] = 1709
         "0011010011101" when "1010011", -- t[83] = 1693
         "0011010001110" when "1010100", -- t[84] = 1678
         "0011001111111" when "1010101", -- t[85] = 1663
         "0011001110000" when "1010110", -- t[86] = 1648
         "0011001100001" when "1010111", -- t[87] = 1633
         "0011001010011" when "1011000", -- t[88] = 1619
         "0011001000100" when "1011001", -- t[89] = 1604
         "0011000110110" when "1011010", -- t[90] = 1590
         "0011000101001" when "1011011", -- t[91] = 1577
         "0011000011011" when "1011100", -- t[92] = 1563
         "0011000001110" when "1011101", -- t[93] = 1550
         "0011000000000" when "1011110", -- t[94] = 1536
         "0010111110011" when "1011111", -- t[95] = 1523
         "0010111100110" when "1100000", -- t[96] = 1510
         "0010111011010" when "1100001", -- t[97] = 1498
         "0010111001101" when "1100010", -- t[98] = 1485
         "0010111000001" when "1100011", -- t[99] = 1473
         "0010110110101" when "1100100", -- t[100] = 1461
         "0010110101001" when "1100101", -- t[101] = 1449
         "0010110011101" when "1100110", -- t[102] = 1437
         "0010110010001" when "1100111", -- t[103] = 1425
         "0010110000110" when "1101000", -- t[104] = 1414
         "0010101111010" when "1101001", -- t[105] = 1402
         "0010101101111" when "1101010", -- t[106] = 1391
         "0010101100100" when "1101011", -- t[107] = 1380
         "0010101011001" when "1101100", -- t[108] = 1369
         "0010101001110" when "1101101", -- t[109] = 1358
         "0010101000100" when "1101110", -- t[110] = 1348
         "0010100111001" when "1101111", -- t[111] = 1337
         "0010100101111" when "1110000", -- t[112] = 1327
         "0010100100101" when "1110001", -- t[113] = 1317
         "0010100011010" when "1110010", -- t[114] = 1306
         "0010100010000" when "1110011", -- t[115] = 1296
         "0010100000111" when "1110100", -- t[116] = 1287
         "0010011111101" when "1110101", -- t[117] = 1277
         "0010011110011" when "1110110", -- t[118] = 1267
         "0010011101010" when "1110111", -- t[119] = 1258
         "0010011100000" when "1111000", -- t[120] = 1248
         "0010011010111" when "1111001", -- t[121] = 1239
         "0010011001110" when "1111010", -- t[122] = 1230
         "0010011000101" when "1111011", -- t[123] = 1221
         "0010010111100" when "1111100", -- t[124] = 1212
         "0010010110011" when "1111101", -- t[125] = 1203
         "0010010101011" when "1111110", -- t[126] = 1195
         "0010010100010" when "1111111", -- t[127] = 1186
         "-------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 7; beta_1 = 9; lambda_1 = 9;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 7; rho_1,1 = 0; sigma_1,1 = 9; wO_1,1 = 13.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_16_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(8 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_16_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(7 downto 0);
  signal s      : std_logic_vector(8 downto 0);
  component fp_log_log_16_t1_pow is
    port ( x : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(7 downto 0);
  signal k_1    : std_logic_vector(12 downto 0);
  signal r0_1   : std_logic_vector(22 downto 0);
  signal r_1    : std_logic_vector(19 downto 0);
  component fp_log_log_16_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;
begin
  sign <= not b(8);
  b0 <= b(7 downto 0) xor (7 downto 0 => sign);

  pow : fp_log_log_16_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(8);
  s_1 <= s(7 downto 0) xor (7 downto 0 => sign_1);
  t_1 : fp_log_log_16_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(12 downto 0) <=
    r0_1(22 downto 10) xor (22 downto 10 => (not (sign xor sign_1)));
  r_1(19 downto 13) <= (19 downto 13 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- TermROM instance for order-2 term.
-- Decomposition:
--   alpha_2 = 3; beta_2 = 4 (1+3); wO_2 = 4.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_16_t2 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_16_t2 is
  signal sign : std_logic;
  signal b0   : std_logic_vector(2 downto 0);
  signal x0   : std_logic_vector(5 downto 0);
  signal r0   : std_logic_vector(3 downto 0);
begin
  sign <= not b(3);
  b0 <= b(2 downto 0) xor (2 downto 0 => sign);
  x0 <= a & b0;

  with x0 select
    r0 <= "0000" when "000000", -- t[0] = 0
          "0000" when "000001", -- t[1] = 0
          "0001" when "000010", -- t[2] = 1
          "0001" when "000011", -- t[3] = 1
          "0011" when "000100", -- t[4] = 3
          "0100" when "000101", -- t[5] = 4
          "0110" when "000110", -- t[6] = 6
          "1000" when "000111", -- t[7] = 8
          "0000" when "001000", -- t[8] = 0
          "0000" when "001001", -- t[9] = 0
          "0000" when "001010", -- t[10] = 0
          "0001" when "001011", -- t[11] = 1
          "0010" when "001100", -- t[12] = 2
          "0011" when "001101", -- t[13] = 3
          "0100" when "001110", -- t[14] = 4
          "0101" when "001111", -- t[15] = 5
          "0000" when "010000", -- t[16] = 0
          "0000" when "010001", -- t[17] = 0
          "0000" when "010010", -- t[18] = 0
          "0000" when "010011", -- t[19] = 0
          "0001" when "010100", -- t[20] = 1
          "0010" when "010101", -- t[21] = 2
          "0010" when "010110", -- t[22] = 2
          "0011" when "010111", -- t[23] = 3
          "0000" when "011000", -- t[24] = 0
          "0000" when "011001", -- t[25] = 0
          "0000" when "011010", -- t[26] = 0
          "0000" when "011011", -- t[27] = 0
          "0001" when "011100", -- t[28] = 1
          "0001" when "011101", -- t[29] = 1
          "0010" when "011110", -- t[30] = 2
          "0010" when "011111", -- t[31] = 2
          "0000" when "100000", -- t[32] = 0
          "0000" when "100001", -- t[33] = 0
          "0000" when "100010", -- t[34] = 0
          "0000" when "100011", -- t[35] = 0
          "0000" when "100100", -- t[36] = 0
          "0001" when "100101", -- t[37] = 1
          "0001" when "100110", -- t[38] = 1
          "0010" when "100111", -- t[39] = 2
          "0000" when "101000", -- t[40] = 0
          "0000" when "101001", -- t[41] = 0
          "0000" when "101010", -- t[42] = 0
          "0000" when "101011", -- t[43] = 0
          "0000" when "101100", -- t[44] = 0
          "0000" when "101101", -- t[45] = 0
          "0001" when "101110", -- t[46] = 1
          "0001" when "101111", -- t[47] = 1
          "0000" when "110000", -- t[48] = 0
          "0000" when "110001", -- t[49] = 0
          "0000" when "110010", -- t[50] = 0
          "0000" when "110011", -- t[51] = 0
          "0000" when "110100", -- t[52] = 0
          "0000" when "110101", -- t[53] = 0
          "0000" when "110110", -- t[54] = 0
          "0001" when "110111", -- t[55] = 1
          "0000" when "111000", -- t[56] = 0
          "0000" when "111001", -- t[57] = 0
          "0000" when "111010", -- t[58] = 0
          "0000" when "111011", -- t[59] = 0
          "0000" when "111100", -- t[60] = 0
          "0000" when "111101", -- t[61] = 0
          "0000" when "111110", -- t[62] = 0
          "0001" when "111111", -- t[63] = 1
          "----" when others;

  r(3 downto 0) <= r0;
  r(19 downto 4) <= (19 downto 4 => ('0'));
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_16 is
  port ( x : in  std_logic_vector(15 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_16 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(19 downto 0);
  component fp_log_log_16_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

  signal a_1 : std_logic_vector(6 downto 0);
  signal b_1 : std_logic_vector(8 downto 0);
  signal r_1 : std_logic_vector(19 downto 0);
  component fp_log_log_16_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(8 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

  signal a_2 : std_logic_vector(2 downto 0);
  signal b_2 : std_logic_vector(3 downto 0);
  signal r_2 : std_logic_vector(19 downto 0);
  component fp_log_log_16_t2 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;

begin
  a_0 <= x(15 downto 9);
  t_0 : fp_log_log_16_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(15 downto 9);
  b_1 <= x(8 downto 0);
  t_1 : fp_log_log_16_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(15 downto 13);
  b_2 <= x(8 downto 5);
  t_2 : fp_log_log_16_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 17; wO = 17.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 10;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 7; beta_1 = 10;
--   T_2 (PowMult): alpha_2 = 4; beta_2 = 5.
-- Guard bits: g = 3.
-- Command line: logfp 17 17 2   rom 7 0   pm 7 10  ah 10 10 10  1 0  7 10 0   pm 4 5  ah 5 10 6  1 1  4 3 0  1 3 3


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 21.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(20 downto 0) );
end entity;

architecture arch of fp_log_log_17_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(20 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "101100001101011000000" when "0000000", -- t[0] = 1448640
          "101011111010000111011" when "0000001", -- t[1] = 1438779
          "101011100111001110010" when "0000010", -- t[2] = 1429106
          "101011010100101011110" when "0000011", -- t[3] = 1419614
          "101011000010011111011" when "0000100", -- t[4] = 1410299
          "101010110000101000010" when "0000101", -- t[5] = 1401154
          "101010011111000101111" when "0000110", -- t[6] = 1392175
          "101010001101110111100" when "0000111", -- t[7] = 1383356
          "101001111100111101000" when "0001000", -- t[8] = 1374696
          "101001101100010100111" when "0001001", -- t[9] = 1366183
          "101001011011111111000" when "0001010", -- t[10] = 1357816
          "101001001011111010111" when "0001011", -- t[11] = 1349591
          "101000111100000111111" when "0001100", -- t[12] = 1341503
          "101000101100100101110" when "0001101", -- t[13] = 1333550
          "101000011101010011111" when "0001110", -- t[14] = 1325727
          "101000001110010001111" when "0001111", -- t[15] = 1318031
          "100111111111011111100" when "0010000", -- t[16] = 1310460
          "100111110000111011111" when "0010001", -- t[17] = 1303007
          "100111100010100110110" when "0010010", -- t[18] = 1295670
          "100111010100011111110" when "0010011", -- t[19] = 1288446
          "100111000110100110101" when "0010100", -- t[20] = 1281333
          "100110111000111010111" when "0010101", -- t[21] = 1274327
          "100110101011011100010" when "0010110", -- t[22] = 1267426
          "100110011110001010100" when "0010111", -- t[23] = 1260628
          "100110010001000101011" when "0011000", -- t[24] = 1253931
          "100110000100001100001" when "0011001", -- t[25] = 1247329
          "100101110111011110110" when "0011010", -- t[26] = 1240822
          "100101101010111101000" when "0011011", -- t[27] = 1234408
          "100101011110100110100" when "0011100", -- t[28] = 1228084
          "100101010010011011000" when "0011101", -- t[29] = 1221848
          "100101000110011010010" when "0011110", -- t[30] = 1215698
          "100100111010100100000" when "0011111", -- t[31] = 1209632
          "100100101110111000001" when "0100000", -- t[32] = 1203649
          "100100100011010110010" when "0100001", -- t[33] = 1197746
          "100100010111111110000" when "0100010", -- t[34] = 1191920
          "100100001100101111100" when "0100011", -- t[35] = 1186172
          "100100000001101010010" when "0100100", -- t[36] = 1180498
          "100011110110101110010" when "0100101", -- t[37] = 1174898
          "100011101011111011001" when "0100110", -- t[38] = 1169369
          "100011100001010000110" when "0100111", -- t[39] = 1163910
          "100011010110101111010" when "0101000", -- t[40] = 1158522
          "100011001100010101111" when "0101001", -- t[41] = 1153199
          "100011000010000100110" when "0101010", -- t[42] = 1147942
          "100010110111111011110" when "0101011", -- t[43] = 1142750
          "100010101101111010100" when "0101100", -- t[44] = 1137620
          "100010100100000001001" when "0101101", -- t[45] = 1132553
          "100010011010001111010" when "0101110", -- t[46] = 1127546
          "100010010000100100110" when "0101111", -- t[47] = 1122598
          "100010000111000001101" when "0110000", -- t[48] = 1117709
          "100001111101100101101" when "0110001", -- t[49] = 1112877
          "100001110100010000100" when "0110010", -- t[50] = 1108100
          "100001101011000010010" when "0110011", -- t[51] = 1103378
          "100001100001111010110" when "0110100", -- t[52] = 1098710
          "100001011000111001110" when "0110101", -- t[53] = 1094094
          "100001001111111111011" when "0110110", -- t[54] = 1089531
          "100001000111001011010" when "0110111", -- t[55] = 1085018
          "100000111110011101011" when "0111000", -- t[56] = 1080555
          "100000110101110101101" when "0111001", -- t[57] = 1076141
          "100000101101010011111" when "0111010", -- t[58] = 1071775
          "100000100100110111111" when "0111011", -- t[59] = 1067455
          "100000011100100001110" when "0111100", -- t[60] = 1063182
          "100000010100010001011" when "0111101", -- t[61] = 1058955
          "100000001100000110100" when "0111110", -- t[62] = 1054772
          "100000000100000001001" when "0111111", -- t[63] = 1050633
          "011111111100000001001" when "1000000", -- t[64] = 1046537
          "011111110100000110011" when "1000001", -- t[65] = 1042483
          "011111101100010000111" when "1000010", -- t[66] = 1038471
          "011111100100100000100" when "1000011", -- t[67] = 1034500
          "011111011100110101000" when "1000100", -- t[68] = 1030568
          "011111010101001110100" when "1000101", -- t[69] = 1026676
          "011111001101101101000" when "1000110", -- t[70] = 1022824
          "011111000110010000001" when "1000111", -- t[71] = 1019009
          "011110111110111000000" when "1001000", -- t[72] = 1015232
          "011110110111100100100" when "1001001", -- t[73] = 1011492
          "011110110000010101100" when "1001010", -- t[74] = 1007788
          "011110101001001010111" when "1001011", -- t[75] = 1004119
          "011110100010000100110" when "1001100", -- t[76] = 1000486
          "011110011011000010111" when "1001101", -- t[77] = 996887
          "011110010100000101011" when "1001110", -- t[78] = 993323
          "011110001101001100000" when "1001111", -- t[79] = 989792
          "011110000110010110110" when "1010000", -- t[80] = 986294
          "011101111111100101101" when "1010001", -- t[81] = 982829
          "011101111000111000011" when "1010010", -- t[82] = 979395
          "011101110010001111001" when "1010011", -- t[83] = 975993
          "011101101011101001101" when "1010100", -- t[84] = 972621
          "011101100101001000001" when "1010101", -- t[85] = 969281
          "011101011110101010010" when "1010110", -- t[86] = 965970
          "011101011000010000001" when "1010111", -- t[87] = 962689
          "011101010001111001101" when "1011000", -- t[88] = 959437
          "011101001011100110110" when "1011001", -- t[89] = 956214
          "011101000101010111011" when "1011010", -- t[90] = 953019
          "011100111111001011100" when "1011011", -- t[91] = 949852
          "011100111001000011000" when "1011100", -- t[92] = 946712
          "011100110010111110000" when "1011101", -- t[93] = 943600
          "011100101100111100010" when "1011110", -- t[94] = 940514
          "011100100110111101111" when "1011111", -- t[95] = 937455
          "011100100001000010101" when "1100000", -- t[96] = 934421
          "011100011011001010110" when "1100001", -- t[97] = 931414
          "011100010101010101111" when "1100010", -- t[98] = 928431
          "011100001111100100001" when "1100011", -- t[99] = 925473
          "011100001001110101011" when "1100100", -- t[100] = 922539
          "011100000100001001110" when "1100101", -- t[101] = 919630
          "011011111110100001001" when "1100110", -- t[102] = 916745
          "011011111000111011011" when "1100111", -- t[103] = 913883
          "011011110011011000101" when "1101000", -- t[104] = 911045
          "011011101101111000101" when "1101001", -- t[105] = 908229
          "011011101000011011100" when "1101010", -- t[106] = 905436
          "011011100011000001001" when "1101011", -- t[107] = 902665
          "011011011101101001100" when "1101100", -- t[108] = 899916
          "011011011000010100101" when "1101101", -- t[109] = 897189
          "011011010011000010011" when "1101110", -- t[110] = 894483
          "011011001101110010110" when "1101111", -- t[111] = 891798
          "011011001000100101111" when "1110000", -- t[112] = 889135
          "011011000011011011100" when "1110001", -- t[113] = 886492
          "011010111110010011101" when "1110010", -- t[114] = 883869
          "011010111001001110010" when "1110011", -- t[115] = 881266
          "011010110100001011011" when "1110100", -- t[116] = 878683
          "011010101111001010111" when "1110101", -- t[117] = 876119
          "011010101010001100111" when "1110110", -- t[118] = 873575
          "011010100101010001010" when "1110111", -- t[119] = 871050
          "011010100000011000000" when "1111000", -- t[120] = 868544
          "011010011011100001000" when "1111001", -- t[121] = 866056
          "011010010110101100011" when "1111010", -- t[122] = 863587
          "011010010001111010000" when "1111011", -- t[123] = 861136
          "011010001101001001111" when "1111100", -- t[124] = 858703
          "011010001000011011111" when "1111101", -- t[125] = 856287
          "011010000011110000001" when "1111110", -- t[126] = 853889
          "011001111111000110100" when "1111111", -- t[127] = 851508
          "---------------------" when others;

  r(20 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 10; mu_1 = 10; lambda_1 = 10.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t1_pow is
  port ( x : in  std_logic_vector(8 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of fp_log_log_17_t1_pow is
  signal pp0 : std_logic_vector(8 downto 0);
  signal r0 : std_logic_vector(8 downto 0);
begin
  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(8 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 7; wO_1,1 = 14.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t1_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_17_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "10011011100101" when "0000000", -- t[0] = 9957
         "10011000100110" when "0000001", -- t[1] = 9766
         "10010101101101" when "0000010", -- t[2] = 9581
         "10010010111010" when "0000011", -- t[3] = 9402
         "10010000001101" when "0000100", -- t[4] = 9229
         "10001101100101" when "0000101", -- t[5] = 9061
         "10001011000010" when "0000110", -- t[6] = 8898
         "10001000100100" when "0000111", -- t[7] = 8740
         "10000110001011" when "0001000", -- t[8] = 8587
         "10000011110111" when "0001001", -- t[9] = 8439
         "10000001100111" when "0001010", -- t[10] = 8295
         "01111111011011" when "0001011", -- t[11] = 8155
         "01111101010011" when "0001100", -- t[12] = 8019
         "01111011001111" when "0001101", -- t[13] = 7887
         "01111001001111" when "0001110", -- t[14] = 7759
         "01110111010010" when "0001111", -- t[15] = 7634
         "01110101011001" when "0010000", -- t[16] = 7513
         "01110011100011" when "0010001", -- t[17] = 7395
         "01110001110000" when "0010010", -- t[18] = 7280
         "01110000000000" when "0010011", -- t[19] = 7168
         "01101110010011" when "0010100", -- t[20] = 7059
         "01101100101000" when "0010101", -- t[21] = 6952
         "01101011000001" when "0010110", -- t[22] = 6849
         "01101001011100" when "0010111", -- t[23] = 6748
         "01100111111010" when "0011000", -- t[24] = 6650
         "01100110011010" when "0011001", -- t[25] = 6554
         "01100100111100" when "0011010", -- t[26] = 6460
         "01100011100001" when "0011011", -- t[27] = 6369
         "01100010001000" when "0011100", -- t[28] = 6280
         "01100000110001" when "0011101", -- t[29] = 6193
         "01011111011100" when "0011110", -- t[30] = 6108
         "01011110001001" when "0011111", -- t[31] = 6025
         "01011100110111" when "0100000", -- t[32] = 5943
         "01011011101000" when "0100001", -- t[33] = 5864
         "01011010011011" when "0100010", -- t[34] = 5787
         "01011001001111" when "0100011", -- t[35] = 5711
         "01011000000101" when "0100100", -- t[36] = 5637
         "01010110111100" when "0100101", -- t[37] = 5564
         "01010101110101" when "0100110", -- t[38] = 5493
         "01010100110000" when "0100111", -- t[39] = 5424
         "01010011101100" when "0101000", -- t[40] = 5356
         "01010010101001" when "0101001", -- t[41] = 5289
         "01010001101000" when "0101010", -- t[42] = 5224
         "01010000101001" when "0101011", -- t[43] = 5161
         "01001111101010" when "0101100", -- t[44] = 5098
         "01001110101101" when "0101101", -- t[45] = 5037
         "01001101110001" when "0101110", -- t[46] = 4977
         "01001100110110" when "0101111", -- t[47] = 4918
         "01001011111101" when "0110000", -- t[48] = 4861
         "01001011000100" when "0110001", -- t[49] = 4804
         "01001010001101" when "0110010", -- t[50] = 4749
         "01001001010111" when "0110011", -- t[51] = 4695
         "01001000100010" when "0110100", -- t[52] = 4642
         "01000111101101" when "0110101", -- t[53] = 4589
         "01000110111010" when "0110110", -- t[54] = 4538
         "01000110001000" when "0110111", -- t[55] = 4488
         "01000101010111" when "0111000", -- t[56] = 4439
         "01000100100110" when "0111001", -- t[57] = 4390
         "01000011110111" when "0111010", -- t[58] = 4343
         "01000011001000" when "0111011", -- t[59] = 4296
         "01000010011010" when "0111100", -- t[60] = 4250
         "01000001101101" when "0111101", -- t[61] = 4205
         "01000001000001" when "0111110", -- t[62] = 4161
         "01000000010101" when "0111111", -- t[63] = 4117
         "00111111101011" when "1000000", -- t[64] = 4075
         "00111111000001" when "1000001", -- t[65] = 4033
         "00111110011000" when "1000010", -- t[66] = 3992
         "00111101101111" when "1000011", -- t[67] = 3951
         "00111101000111" when "1000100", -- t[68] = 3911
         "00111100100000" when "1000101", -- t[69] = 3872
         "00111011111010" when "1000110", -- t[70] = 3834
         "00111011010100" when "1000111", -- t[71] = 3796
         "00111010101111" when "1001000", -- t[72] = 3759
         "00111010001010" when "1001001", -- t[73] = 3722
         "00111001100110" when "1001010", -- t[74] = 3686
         "00111001000011" when "1001011", -- t[75] = 3651
         "00111000100000" when "1001100", -- t[76] = 3616
         "00110111111101" when "1001101", -- t[77] = 3581
         "00110111011100" when "1001110", -- t[78] = 3548
         "00110110111010" when "1001111", -- t[79] = 3514
         "00110110011010" when "1010000", -- t[80] = 3482
         "00110101111010" when "1010001", -- t[81] = 3450
         "00110101011010" when "1010010", -- t[82] = 3418
         "00110100111011" when "1010011", -- t[83] = 3387
         "00110100011100" when "1010100", -- t[84] = 3356
         "00110011111110" when "1010101", -- t[85] = 3326
         "00110011100000" when "1010110", -- t[86] = 3296
         "00110011000010" when "1010111", -- t[87] = 3266
         "00110010100101" when "1011000", -- t[88] = 3237
         "00110010001001" when "1011001", -- t[89] = 3209
         "00110001101101" when "1011010", -- t[90] = 3181
         "00110001010001" when "1011011", -- t[91] = 3153
         "00110000110110" when "1011100", -- t[92] = 3126
         "00110000011011" when "1011101", -- t[93] = 3099
         "00110000000001" when "1011110", -- t[94] = 3073
         "00101111100110" when "1011111", -- t[95] = 3046
         "00101111001101" when "1100000", -- t[96] = 3021
         "00101110110011" when "1100001", -- t[97] = 2995
         "00101110011010" when "1100010", -- t[98] = 2970
         "00101110000010" when "1100011", -- t[99] = 2946
         "00101101101001" when "1100100", -- t[100] = 2921
         "00101101010001" when "1100101", -- t[101] = 2897
         "00101100111010" when "1100110", -- t[102] = 2874
         "00101100100010" when "1100111", -- t[103] = 2850
         "00101100001011" when "1101000", -- t[104] = 2827
         "00101011110100" when "1101001", -- t[105] = 2804
         "00101011011110" when "1101010", -- t[106] = 2782
         "00101011001000" when "1101011", -- t[107] = 2760
         "00101010110010" when "1101100", -- t[108] = 2738
         "00101010011100" when "1101101", -- t[109] = 2716
         "00101010000111" when "1101110", -- t[110] = 2695
         "00101001110010" when "1101111", -- t[111] = 2674
         "00101001011101" when "1110000", -- t[112] = 2653
         "00101001001001" when "1110001", -- t[113] = 2633
         "00101000110101" when "1110010", -- t[114] = 2613
         "00101000100001" when "1110011", -- t[115] = 2593
         "00101000001101" when "1110100", -- t[116] = 2573
         "00100111111010" when "1110101", -- t[117] = 2554
         "00100111100111" when "1110110", -- t[118] = 2535
         "00100111010100" when "1110111", -- t[119] = 2516
         "00100111000001" when "1111000", -- t[120] = 2497
         "00100110101110" when "1111001", -- t[121] = 2478
         "00100110011100" when "1111010", -- t[122] = 2460
         "00100110001010" when "1111011", -- t[123] = 2442
         "00100101111000" when "1111100", -- t[124] = 2424
         "00100101100111" when "1111101", -- t[125] = 2407
         "00100101010101" when "1111110", -- t[126] = 2389
         "00100101000100" when "1111111", -- t[127] = 2372
         "--------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 7; beta_1 = 10; lambda_1 = 10;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 7; rho_1,1 = 0; sigma_1,1 = 10; wO_1,1 = 14.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(9 downto 0);
         r : out std_logic_vector(20 downto 0) );
end entity;

architecture arch of fp_log_log_17_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(8 downto 0);
  signal s      : std_logic_vector(9 downto 0);
  component fp_log_log_17_t1_pow is
    port ( x : in  std_logic_vector(8 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(8 downto 0);
  signal k_1    : std_logic_vector(13 downto 0);
  signal r0_1   : std_logic_vector(24 downto 0);
  signal r_1    : std_logic_vector(20 downto 0);
  component fp_log_log_17_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;
begin
  sign <= not b(9);
  b0 <= b(8 downto 0) xor (8 downto 0 => sign);

  pow : fp_log_log_17_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(9);
  s_1 <= s(8 downto 0) xor (8 downto 0 => sign_1);
  t_1 : fp_log_log_17_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(13 downto 0) <=
    r0_1(24 downto 11) xor (24 downto 11 => (not (sign xor sign_1)));
  r_1(20 downto 14) <= (20 downto 14 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 5; mu_2 = 10; lambda_2 = 6.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t2_pow is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_log_log_17_t2_pow is
  signal pp0 : std_logic_vector(8 downto 0);
  signal pp1 : std_logic_vector(8 downto 0);
  signal pp2 : std_logic_vector(8 downto 0);
  signal r0 : std_logic_vector(8 downto 0);
begin
  pp0(8) <= '0';
  pp1(8) <= '0';
  pp2(8) <= '0';

  pp0(7) <= x(2) and x(3);
  pp1(7) <= x(3);
  pp2(7) <= '0';

  pp0(6) <= x(1) and x(3);
  pp1(6) <= '0';
  pp2(6) <= '0';

  pp0(5) <= x(0) and x(3);
  pp1(5) <= x(1) and x(2);
  pp2(5) <= x(2);

  pp0(4) <= x(0) and x(2);
  pp1(4) <= x(3);
  pp2(4) <= '0';

  pp0(3) <= x(0) and x(1);
  pp1(3) <= x(1);
  pp2(3) <= x(2);

  pp0(2) <= x(0);
  pp1(2) <= x(1);
  pp2(2) <= '0';

  pp0(1) <= '0';
  pp1(1) <= '0';
  pp2(1) <= '0';

  pp0(0) <= '0';
  pp1(0) <= '0';
  pp2(0) <= '0';

  r0 <= pp0 + pp1 + pp2;
  r <= "1" & r0(8 downto 4);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 4; wO_2,1 = 6.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t2_t1 is
  port ( a : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of fp_log_log_17_t2_t1 is
  signal x : std_logic_vector(3 downto 0);
begin
  x <= a;

  with x select
    r <= "101100" when "0000", -- t[0] = 44
         "100010" when "0001", -- t[1] = 34
         "011011" when "0010", -- t[2] = 27
         "010110" when "0011", -- t[3] = 22
         "010011" when "0100", -- t[4] = 19
         "010000" when "0101", -- t[5] = 16
         "001101" when "0110", -- t[6] = 13
         "001011" when "0111", -- t[7] = 11
         "001010" when "1000", -- t[8] = 10
         "001001" when "1001", -- t[9] = 9
         "001000" when "1010", -- t[10] = 8
         "000111" when "1011", -- t[11] = 7
         "000110" when "1100", -- t[12] = 6
         "000101" when "1101", -- t[13] = 5
         "000101" when "1110", -- t[14] = 5
         "000100" when "1111", -- t[15] = 4
         "------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_2.
-- Decomposition:
--   alpha_2,2 = 1; sigma'_2,2 = 2; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t2_t2 is
  port ( a : in  std_logic_vector(0 downto 0);
         s : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of fp_log_log_17_t2_t2 is
  signal x : std_logic_vector(2 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0" when "000", -- t[0] = 0
         "0" when "001", -- t[1] = 0
         "1" when "010", -- t[2] = 1
         "1" when "011", -- t[3] = 1
         "0" when "100", -- t[4] = 0
         "0" when "101", -- t[5] = 0
         "0" when "110", -- t[6] = 0
         "0" when "111", -- t[7] = 0
         "-" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 4; beta_2 = 5; lambda_2 = 6;  m_2 = 2;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 4; rho_2,1 = 0; sigma_2,1 = 3; wO_2,1 = 6;
--   Q_2,2 (ROM):  alpha_2,2 = 1; rho_2,2 = 3; sigma_2,2 = 3; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17_t2 is
  port ( a : in  std_logic_vector(3 downto 0);
         b : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(20 downto 0) );
end entity;

architecture arch of fp_log_log_17_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(3 downto 0);
  signal s      : std_logic_vector(5 downto 0);
  component fp_log_log_17_t2_pow is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  signal a_1    : std_logic_vector(3 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(1 downto 0);
  signal k_1    : std_logic_vector(5 downto 0);
  signal r0_1   : std_logic_vector(9 downto 0);
  signal r_1    : std_logic_vector(20 downto 0);
  component fp_log_log_17_t2_t1 is
    port ( a : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  signal a_2    : std_logic_vector(0 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(1 downto 0);
  signal r0_2   : std_logic_vector(0 downto 0);
  signal r_2    : std_logic_vector(20 downto 0);
  component fp_log_log_17_t2_t2 is
    port ( a : in  std_logic_vector(0 downto 0);
           s : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;
begin
  sign <= not b(4);
  b0 <= b(3 downto 0) xor (3 downto 0 => sign);

  pow : fp_log_log_17_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(3 downto 0);
  sign_1 <= not s(5);
  s_1 <= s(4 downto 3) xor (4 downto 3 => sign_1);
  t_1 : fp_log_log_17_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(5 downto 0) <=
    r0_1(9 downto 4) xor (9 downto 4 => ((sign_1)));
  r_1(20 downto 6) <= (20 downto 6 => ((sign_1)));

  a_2 <= a(3 downto 3);
  sign_2 <= not s(2);
  s_2 <= s(1 downto 0) xor (1 downto 0 => sign_2);
  t_2 : fp_log_log_17_t2_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(0 downto 0) <=
    r0_2 xor (0 downto 0 => ((sign_2)));
  r_2(20 downto 1) <= (20 downto 1 => ((sign_2)));

  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_17 is
  port ( x : in  std_logic_vector(16 downto 0);
         r : out std_logic_vector(20 downto 0) );
end entity;

architecture arch of fp_log_log_17 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(20 downto 0);
  component fp_log_log_17_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(20 downto 0) );
  end component;

  signal a_1 : std_logic_vector(6 downto 0);
  signal b_1 : std_logic_vector(9 downto 0);
  signal r_1 : std_logic_vector(20 downto 0);
  component fp_log_log_17_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(20 downto 0) );
  end component;

  signal a_2 : std_logic_vector(3 downto 0);
  signal b_2 : std_logic_vector(4 downto 0);
  signal r_2 : std_logic_vector(20 downto 0);
  component fp_log_log_17_t2 is
    port ( a : in  std_logic_vector(3 downto 0);
           b : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(20 downto 0) );
  end component;

begin
  a_0 <= x(16 downto 10);
  t_0 : fp_log_log_17_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(16 downto 10);
  b_1 <= x(9 downto 0);
  t_1 : fp_log_log_17_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(16 downto 13);
  b_2 <= x(9 downto 5);
  t_2 : fp_log_log_17_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 18; wO = 18.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 11;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 7; beta_1 = 11;
--   T_2 (PowMult): alpha_2 = 5; beta_2 = 6.
-- Guard bits: g = 3.
-- Command line: logfp 18 18 2   rom 7 0   pm 7 11  ah 11 11 11  1 0  7 11 0   pm 5 6  ah 6 12 10  1 1  5 6 0  2 4 6


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 22.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(21 downto 0) );
end entity;

architecture arch of fp_log_log_18_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(21 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "1011000011010101111000" when "0000000", -- t[0] = 2897272
          "1010111110100001101110" when "0000001", -- t[1] = 2877550
          "1010111001110011011011" when "0000010", -- t[2] = 2858203
          "1010110101001010110100" when "0000011", -- t[3] = 2839220
          "1010110000100111110010" when "0000100", -- t[4] = 2820594
          "1010101100001010000001" when "0000101", -- t[5] = 2802305
          "1010100111110001011010" when "0000110", -- t[6] = 2784346
          "1010100011011101110100" when "0000111", -- t[7] = 2766708
          "1010011111001111001000" when "0001000", -- t[8] = 2749384
          "1010011011000101000110" when "0001001", -- t[9] = 2732358
          "1010010110111111101000" when "0001010", -- t[10] = 2715624
          "1010010010111110100110" when "0001011", -- t[11] = 2699174
          "1010001111000001111011" when "0001100", -- t[12] = 2683003
          "1010001011001001011001" when "0001101", -- t[13] = 2667097
          "1010000111010100111011" when "0001110", -- t[14] = 2651451
          "1010000011100100011010" when "0001111", -- t[15] = 2636058
          "1001111111110111110010" when "0010000", -- t[16] = 2620914
          "1001111100001110110111" when "0010001", -- t[17] = 2606007
          "1001111000101001100101" when "0010010", -- t[18] = 2591333
          "1001110101000111110110" when "0010011", -- t[19] = 2576886
          "1001110001101001100110" when "0010100", -- t[20] = 2562662
          "1001101110001110101011" when "0010101", -- t[21] = 2548651
          "1001101010110111000001" when "0010110", -- t[22] = 2534849
          "1001100111100010100100" when "0010111", -- t[23] = 2521252
          "1001100100010001010001" when "0011000", -- t[24] = 2507857
          "1001100001000010111101" when "0011001", -- t[25] = 2494653
          "1001011101110111100111" when "0011010", -- t[26] = 2481639
          "1001011010101111001011" when "0011011", -- t[27] = 2468811
          "1001010111101001100100" when "0011100", -- t[28] = 2456164
          "1001010100100110101100" when "0011101", -- t[29] = 2443692
          "1001010001100110100000" when "0011110", -- t[30] = 2431392
          "1001001110101000111100" when "0011111", -- t[31] = 2419260
          "1001001011101101111110" when "0100000", -- t[32] = 2407294
          "1001001000110101011110" when "0100001", -- t[33] = 2395486
          "1001000101111111011100" when "0100010", -- t[34] = 2383836
          "1001000011001011110011" when "0100011", -- t[35] = 2372339
          "1001000000011010100001" when "0100100", -- t[36] = 2360993
          "1000111101101011100000" when "0100101", -- t[37] = 2349792
          "1000111010111110101110" when "0100110", -- t[38] = 2338734
          "1000111000010100001001" when "0100111", -- t[39] = 2327817
          "1000110101101011101111" when "0101000", -- t[40] = 2317039
          "1000110011000101011001" when "0101001", -- t[41] = 2306393
          "1000110000100001001000" when "0101010", -- t[42] = 2295880
          "1000101101111110110111" when "0101011", -- t[43] = 2285495
          "1000101011011110100101" when "0101100", -- t[44] = 2275237
          "1000101001000000001110" when "0101101", -- t[45] = 2265102
          "1000100110100011110000" when "0101110", -- t[46] = 2255088
          "1000100100001001001000" when "0101111", -- t[47] = 2245192
          "1000100001110000010110" when "0110000", -- t[48] = 2235414
          "1000011111011001010101" when "0110001", -- t[49] = 2225749
          "1000011101000100000100" when "0110010", -- t[50] = 2216196
          "1000011010110000100000" when "0110011", -- t[51] = 2206752
          "1000011000011110101001" when "0110100", -- t[52] = 2197417
          "1000010110001110011010" when "0110101", -- t[53] = 2188186
          "1000010011111111110010" when "0110110", -- t[54] = 2179058
          "1000010001110010110000" when "0110111", -- t[55] = 2170032
          "1000001111100111010011" when "0111000", -- t[56] = 2161107
          "1000001101011101010110" when "0111001", -- t[57] = 2152278
          "1000001011010100111001" when "0111010", -- t[58] = 2143545
          "1000001001001101111011" when "0111011", -- t[59] = 2134907
          "1000000111001000011001" when "0111100", -- t[60] = 2126361
          "1000000101000100010010" when "0111101", -- t[61] = 2117906
          "1000000011000001100100" when "0111110", -- t[62] = 2109540
          "1000000001000000001110" when "0111111", -- t[63] = 2101262
          "0111111111000000001110" when "1000000", -- t[64] = 2093070
          "0111111101000001100011" when "1000001", -- t[65] = 2084963
          "0111111011000100001010" when "1000010", -- t[66] = 2076938
          "0111111001001000000011" when "1000011", -- t[67] = 2068995
          "0111110111001101001101" when "1000100", -- t[68] = 2061133
          "0111110101010011100110" when "1000101", -- t[69] = 2053350
          "0111110011011011001100" when "1000110", -- t[70] = 2045644
          "0111110001100011111110" when "1000111", -- t[71] = 2038014
          "0111101111101101111100" when "1001000", -- t[72] = 2030460
          "0111101101111001000100" when "1001001", -- t[73] = 2022980
          "0111101100000101010100" when "1001010", -- t[74] = 2015572
          "0111101010010010101011" when "1001011", -- t[75] = 2008235
          "0111101000100001001001" when "1001100", -- t[76] = 2000969
          "0111100110110000101100" when "1001101", -- t[77] = 1993772
          "0111100101000001010011" when "1001110", -- t[78] = 1986643
          "0111100011010010111101" when "1001111", -- t[79] = 1979581
          "0111100001100101101001" when "1010000", -- t[80] = 1972585
          "0111011111111001010110" when "1010001", -- t[81] = 1965654
          "0111011110001110000010" when "1010010", -- t[82] = 1958786
          "0111011100100011101110" when "1010011", -- t[83] = 1951982
          "0111011010111010011000" when "1010100", -- t[84] = 1945240
          "0111011001010001111110" when "1010101", -- t[85] = 1938558
          "0111010111101010100001" when "1010110", -- t[86] = 1931937
          "0111010110000011111111" when "1010111", -- t[87] = 1925375
          "0111010100011110010111" when "1011000", -- t[88] = 1918871
          "0111010010111001101001" when "1011001", -- t[89] = 1912425
          "0111010001010101110011" when "1011010", -- t[90] = 1906035
          "0111001111110010110101" when "1011011", -- t[91] = 1899701
          "0111001110010000101110" when "1011100", -- t[92] = 1893422
          "0111001100101111011101" when "1011101", -- t[93] = 1887197
          "0111001011001111000010" when "1011110", -- t[94] = 1881026
          "0111001001101111011011" when "1011111", -- t[95] = 1874907
          "0111001000010000101000" when "1100000", -- t[96] = 1868840
          "0111000110110010101000" when "1100001", -- t[97] = 1862824
          "0111000101010101011010" when "1100010", -- t[98] = 1856858
          "0111000011111000111111" when "1100011", -- t[99] = 1850943
          "0111000010011101010100" when "1100100", -- t[100] = 1845076
          "0111000001000010011010" when "1100101", -- t[101] = 1839258
          "0110111111101000001111" when "1100110", -- t[102] = 1833487
          "0110111110001110110011" when "1100111", -- t[103] = 1827763
          "0110111100110110000110" when "1101000", -- t[104] = 1822086
          "0110111011011110000111" when "1101001", -- t[105] = 1816455
          "0110111010000110110101" when "1101010", -- t[106] = 1810869
          "0110111000110000001111" when "1101011", -- t[107] = 1805327
          "0110110111011010010101" when "1101100", -- t[108] = 1799829
          "0110110110000101000111" when "1101101", -- t[109] = 1794375
          "0110110100110000100011" when "1101110", -- t[110] = 1788963
          "0110110011011100101010" when "1101111", -- t[111] = 1783594
          "0110110010001001011011" when "1110000", -- t[112] = 1778267
          "0110110000110110110100" when "1110001", -- t[113] = 1772980
          "0110101111100100110110" when "1110010", -- t[114] = 1767734
          "0110101110010011100001" when "1110011", -- t[115] = 1762529
          "0110101101000010110011" when "1110100", -- t[116] = 1757363
          "0110101011110010101100" when "1110101", -- t[117] = 1752236
          "0110101010100011001100" when "1110110", -- t[118] = 1747148
          "0110101001010100010001" when "1110111", -- t[119] = 1742097
          "0110101000000101111101" when "1111000", -- t[120] = 1737085
          "0110100110111000001110" when "1111001", -- t[121] = 1732110
          "0110100101101011000011" when "1111010", -- t[122] = 1727171
          "0110100100011110011101" when "1111011", -- t[123] = 1722269
          "0110100011010010011011" when "1111100", -- t[124] = 1717403
          "0110100010000110111100" when "1111101", -- t[125] = 1712572
          "0110100000111100000000" when "1111110", -- t[126] = 1707776
          "0110011111110001100110" when "1111111", -- t[127] = 1703014
          "----------------------" when others;

  r(21 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 11; mu_1 = 11; lambda_1 = 11.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t1_pow is
  port ( x : in  std_logic_vector(9 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of fp_log_log_18_t1_pow is
  signal pp0 : std_logic_vector(9 downto 0);
  signal r0 : std_logic_vector(9 downto 0);
begin
  pp0(9) <= x(9);

  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(9 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 7; wO_1,1 = 15.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t1_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of fp_log_log_18_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "100110111001010" when "0000000", -- t[0] = 19914
         "100110001001100" when "0000001", -- t[1] = 19532
         "100101011011010" when "0000010", -- t[2] = 19162
         "100100101110100" when "0000011", -- t[3] = 18804
         "100100000011001" when "0000100", -- t[4] = 18457
         "100011011001001" when "0000101", -- t[5] = 18121
         "100010110000100" when "0000110", -- t[6] = 17796
         "100010001001001" when "0000111", -- t[7] = 17481
         "100001100010111" when "0001000", -- t[8] = 17175
         "100000111101110" when "0001001", -- t[9] = 16878
         "100000011001110" when "0001010", -- t[10] = 16590
         "011111110110110" when "0001011", -- t[11] = 16310
         "011111010100110" when "0001100", -- t[12] = 16038
         "011110110011110" when "0001101", -- t[13] = 15774
         "011110010011110" when "0001110", -- t[14] = 15518
         "011101110100100" when "0001111", -- t[15] = 15268
         "011101010110001" when "0010000", -- t[16] = 15025
         "011100111000101" when "0010001", -- t[17] = 14789
         "011100011011111" when "0010010", -- t[18] = 14559
         "011011111111111" when "0010011", -- t[19] = 14335
         "011011100100101" when "0010100", -- t[20] = 14117
         "011011001010001" when "0010101", -- t[21] = 13905
         "011010110000010" when "0010110", -- t[22] = 13698
         "011010010111000" when "0010111", -- t[23] = 13496
         "011001111110011" when "0011000", -- t[24] = 13299
         "011001100110011" when "0011001", -- t[25] = 13107
         "011001001111000" when "0011010", -- t[26] = 12920
         "011000111000010" when "0011011", -- t[27] = 12738
         "011000100001111" when "0011100", -- t[28] = 12559
         "011000001100001" when "0011101", -- t[29] = 12385
         "010111110110111" when "0011110", -- t[30] = 12215
         "010111100010001" when "0011111", -- t[31] = 12049
         "010111001101111" when "0100000", -- t[32] = 11887
         "010110111010000" when "0100001", -- t[33] = 11728
         "010110100110101" when "0100010", -- t[34] = 11573
         "010110010011110" when "0100011", -- t[35] = 11422
         "010110000001001" when "0100100", -- t[36] = 11273
         "010101101111000" when "0100101", -- t[37] = 11128
         "010101011101010" when "0100110", -- t[38] = 10986
         "010101001100000" when "0100111", -- t[39] = 10848
         "010100111011000" when "0101000", -- t[40] = 10712
         "010100101010011" when "0101001", -- t[41] = 10579
         "010100011010001" when "0101010", -- t[42] = 10449
         "010100001010001" when "0101011", -- t[43] = 10321
         "010011111010100" when "0101100", -- t[44] = 10196
         "010011101011010" when "0101101", -- t[45] = 10074
         "010011011100010" when "0101110", -- t[46] = 9954
         "010011001101101" when "0101111", -- t[47] = 9837
         "010010111111010" when "0110000", -- t[48] = 9722
         "010010110001001" when "0110001", -- t[49] = 9609
         "010010100011010" when "0110010", -- t[50] = 9498
         "010010010101110" when "0110011", -- t[51] = 9390
         "010010001000011" when "0110100", -- t[52] = 9283
         "010001111011011" when "0110101", -- t[53] = 9179
         "010001101110100" when "0110110", -- t[54] = 9076
         "010001100010000" when "0110111", -- t[55] = 8976
         "010001010101101" when "0111000", -- t[56] = 8877
         "010001001001100" when "0111001", -- t[57] = 8780
         "010000111101101" when "0111010", -- t[58] = 8685
         "010000110010000" when "0111011", -- t[59] = 8592
         "010000100110100" when "0111100", -- t[60] = 8500
         "010000011011010" when "0111101", -- t[61] = 8410
         "010000010000010" when "0111110", -- t[62] = 8322
         "010000000101011" when "0111111", -- t[63] = 8235
         "001111111010110" when "1000000", -- t[64] = 8150
         "001111110000010" when "1000001", -- t[65] = 8066
         "001111100101111" when "1000010", -- t[66] = 7983
         "001111011011110" when "1000011", -- t[67] = 7902
         "001111010001111" when "1000100", -- t[68] = 7823
         "001111001000000" when "1000101", -- t[69] = 7744
         "001110111110011" when "1000110", -- t[70] = 7667
         "001110110101000" when "1000111", -- t[71] = 7592
         "001110101011101" when "1001000", -- t[72] = 7517
         "001110100010100" when "1001001", -- t[73] = 7444
         "001110011001100" when "1001010", -- t[74] = 7372
         "001110010000101" when "1001011", -- t[75] = 7301
         "001110000111111" when "1001100", -- t[76] = 7231
         "001101111111011" when "1001101", -- t[77] = 7163
         "001101110110111" when "1001110", -- t[78] = 7095
         "001101101110101" when "1001111", -- t[79] = 7029
         "001101100110011" when "1010000", -- t[80] = 6963
         "001101011110011" when "1010001", -- t[81] = 6899
         "001101010110100" when "1010010", -- t[82] = 6836
         "001101001110101" when "1010011", -- t[83] = 6773
         "001101000111000" when "1010100", -- t[84] = 6712
         "001100111111011" when "1010101", -- t[85] = 6651
         "001100111000000" when "1010110", -- t[86] = 6592
         "001100110000101" when "1010111", -- t[87] = 6533
         "001100101001011" when "1011000", -- t[88] = 6475
         "001100100010010" when "1011001", -- t[89] = 6418
         "001100011011010" when "1011010", -- t[90] = 6362
         "001100010100010" when "1011011", -- t[91] = 6306
         "001100001101100" when "1011100", -- t[92] = 6252
         "001100000110110" when "1011101", -- t[93] = 6198
         "001100000000001" when "1011110", -- t[94] = 6145
         "001011111001101" when "1011111", -- t[95] = 6093
         "001011110011001" when "1100000", -- t[96] = 6041
         "001011101100111" when "1100001", -- t[97] = 5991
         "001011100110100" when "1100010", -- t[98] = 5940
         "001011100000011" when "1100011", -- t[99] = 5891
         "001011011010010" when "1100100", -- t[100] = 5842
         "001011010100010" when "1100101", -- t[101] = 5794
         "001011001110011" when "1100110", -- t[102] = 5747
         "001011001000100" when "1100111", -- t[103] = 5700
         "001011000010110" when "1101000", -- t[104] = 5654
         "001010111101001" when "1101001", -- t[105] = 5609
         "001010110111100" when "1101010", -- t[106] = 5564
         "001010110010000" when "1101011", -- t[107] = 5520
         "001010101100100" when "1101100", -- t[108] = 5476
         "001010100111001" when "1101101", -- t[109] = 5433
         "001010100001110" when "1101110", -- t[110] = 5390
         "001010011100100" when "1101111", -- t[111] = 5348
         "001010010111011" when "1110000", -- t[112] = 5307
         "001010010010010" when "1110001", -- t[113] = 5266
         "001010001101010" when "1110010", -- t[114] = 5226
         "001010001000010" when "1110011", -- t[115] = 5186
         "001010000011010" when "1110100", -- t[116] = 5146
         "001001111110100" when "1110101", -- t[117] = 5108
         "001001111001101" when "1110110", -- t[118] = 5069
         "001001110100111" when "1110111", -- t[119] = 5031
         "001001110000010" when "1111000", -- t[120] = 4994
         "001001101011101" when "1111001", -- t[121] = 4957
         "001001100111000" when "1111010", -- t[122] = 4920
         "001001100010100" when "1111011", -- t[123] = 4884
         "001001011110001" when "1111100", -- t[124] = 4849
         "001001011001101" when "1111101", -- t[125] = 4813
         "001001010101011" when "1111110", -- t[126] = 4779
         "001001010001000" when "1111111", -- t[127] = 4744
         "---------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 7; beta_1 = 11; lambda_1 = 11;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 7; rho_1,1 = 0; sigma_1,1 = 11; wO_1,1 = 15.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(21 downto 0) );
end entity;

architecture arch of fp_log_log_18_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(9 downto 0);
  signal s      : std_logic_vector(10 downto 0);
  component fp_log_log_18_t1_pow is
    port ( x : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(9 downto 0);
  signal k_1    : std_logic_vector(14 downto 0);
  signal r0_1   : std_logic_vector(26 downto 0);
  signal r_1    : std_logic_vector(21 downto 0);
  component fp_log_log_18_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(14 downto 0) );
  end component;
begin
  sign <= not b(10);
  b0 <= b(9 downto 0) xor (9 downto 0 => sign);

  pow : fp_log_log_18_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(10);
  s_1 <= s(9 downto 0) xor (9 downto 0 => sign_1);
  t_1 : fp_log_log_18_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(14 downto 0) <=
    r0_1(26 downto 12) xor (26 downto 12 => (not (sign xor sign_1)));
  r_1(21 downto 15) <= (21 downto 15 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_fp_log.all;

entity fp_log_log_18_t1_clk is
  port ( a   : in  std_logic_vector(6 downto 0);
         b   : in  std_logic_vector(10 downto 0);
         r   : out std_logic_vector(21 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_18_t1_clk is
  signal sign_0 : std_logic;
  signal b0_0   : std_logic_vector(9 downto 0);
  signal s_0    : std_logic_vector(10 downto 0);
  component fp_log_log_18_t1_pow is
    port ( x : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  signal a_1_0    : std_logic_vector(6 downto 0);
  signal sign_1_0 : std_logic;
  signal sgn_1_0  : std_logic;
  signal sgn_1_1  : std_logic;
  signal sgn_1_2  : std_logic;
  signal sgn_1_3  : std_logic;
  signal s_1_0    : std_logic_vector(10 downto 0);
  signal s_1_1    : std_logic_vector(10 downto 0);
  signal k_1_0    : std_logic_vector(14 downto 0);
  signal k_1_1    : std_logic_vector(14 downto 0);
  signal r0_1_3   : std_logic_vector(25 downto 0);
  signal r1_1_3   : std_logic_vector(26 downto 0);
  signal r_1_3    : std_logic_vector(21 downto 0);
  component fp_log_log_18_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(14 downto 0) );
  end component;
begin
  sign_0 <= not b(10);
  b0_0 <= b(9 downto 0) xor (9 downto 0 => sign_0);

  pow : fp_log_log_18_t1_pow
    port map ( x => b0_0,
               r => s_0 );

  a_1_0 <= a(6 downto 0);
  sign_1_0 <= not s_0(10);
  sgn_1_0 <= sign_0 xor sign_1_0;
  s_1_0 <= (s_0(9 downto 0) xor (9 downto 0 => sign_1_0)) & "1";
  t_1 : fp_log_log_18_t1_t1
    port map ( a => a_1_0,
               r => k_1_0 );

  mult_r0_1 : mult_clk
    generic map ( wX    => 15,
                  wY    => 11,
                  first => 0,
                  steps => 2 )
    port map ( nX  => k_1_1,
               nY  => s_1_1,
               nR  => r0_1_3,
               clk => clk );
  r1_1_3 <= "0" & r0_1_3;
                 
  r_1_3(14 downto 0) <=
    r1_1_3(26 downto 12) xor (26 downto 12 => (not (sgn_1_3)));
  r_1_3(21 downto 15) <= (21 downto 15 => (not (sgn_1_3)));

  process(clk)
  begin
    if clk'event and clk = '1' then
      s_1_1   <= s_1_0;
      k_1_1   <= k_1_0;
      sgn_1_1 <= sgn_1_0;
      sgn_1_2 <= sgn_1_1;
      sgn_1_3 <= sgn_1_2;
    end if;
  end process;
  
  r <= r_1_3;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 6; mu_2 = 12; lambda_2 = 10.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t2_pow is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of fp_log_log_18_t2_pow is
  signal pp0 : std_logic_vector(10 downto 0);
  signal pp1 : std_logic_vector(10 downto 0);
  signal pp2 : std_logic_vector(10 downto 0);
  signal pp3 : std_logic_vector(10 downto 0);
  signal r0 : std_logic_vector(10 downto 0);
begin
  pp0(10) <= '0';
  pp1(10) <= '0';
  pp2(10) <= '0';
  pp3(10) <= '0';

  pp0(9) <= x(3) and x(4);
  pp1(9) <= x(4);
  pp2(9) <= '0';
  pp3(9) <= '0';

  pp0(8) <= x(2) and x(4);
  pp1(8) <= '0';
  pp2(8) <= '0';
  pp3(8) <= '0';

  pp0(7) <= x(1) and x(4);
  pp1(7) <= x(2) and x(3);
  pp2(7) <= x(3);
  pp3(7) <= '0';

  pp0(6) <= x(0) and x(4);
  pp1(6) <= x(1) and x(3);
  pp2(6) <= '0';
  pp3(6) <= '0';

  pp0(5) <= x(0) and x(3);
  pp1(5) <= x(1) and x(2);
  pp2(5) <= x(2);
  pp3(5) <= x(4);

  pp0(4) <= x(0) and x(2);
  pp1(4) <= x(3);
  pp2(4) <= '0';
  pp3(4) <= '0';

  pp0(3) <= x(0) and x(1);
  pp1(3) <= x(1);
  pp2(3) <= x(2);
  pp3(3) <= '0';

  pp0(2) <= x(0);
  pp1(2) <= x(1);
  pp2(2) <= '0';
  pp3(2) <= '0';

  pp0(1) <= '0';
  pp1(1) <= '0';
  pp2(1) <= '0';
  pp3(1) <= '0';

  pp0(0) <= '0';
  pp1(0) <= '0';
  pp2(0) <= '0';
  pp3(0) <= '0';

  r0 <= pp0 + pp1 + pp2 + pp3;
  r <= "1" & r0(10 downto 2);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 5; wO_2,1 = 7.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t2_t1 is
  port ( a : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_log_log_18_t2_t1 is
  signal x : std_logic_vector(4 downto 0);
begin
  x <= a;

  with x select
    r <= "1011101" when "00000", -- t[0] = 93
         "1010001" when "00001", -- t[1] = 81
         "1001000" when "00010", -- t[2] = 72
         "1000000" when "00011", -- t[3] = 64
         "0111010" when "00100", -- t[4] = 58
         "0110100" when "00101", -- t[5] = 52
         "0101111" when "00110", -- t[6] = 47
         "0101011" when "00111", -- t[7] = 43
         "0100111" when "01000", -- t[8] = 39
         "0100011" when "01001", -- t[9] = 35
         "0100001" when "01010", -- t[10] = 33
         "0011110" when "01011", -- t[11] = 30
         "0011100" when "01100", -- t[12] = 28
         "0011010" when "01101", -- t[13] = 26
         "0011000" when "01110", -- t[14] = 24
         "0010110" when "01111", -- t[15] = 22
         "0010101" when "10000", -- t[16] = 21
         "0010011" when "10001", -- t[17] = 19
         "0010010" when "10010", -- t[18] = 18
         "0010001" when "10011", -- t[19] = 17
         "0010000" when "10100", -- t[20] = 16
         "0001111" when "10101", -- t[21] = 15
         "0001110" when "10110", -- t[22] = 14
         "0001101" when "10111", -- t[23] = 13
         "0001101" when "11000", -- t[24] = 13
         "0001100" when "11001", -- t[25] = 12
         "0001011" when "11010", -- t[26] = 11
         "0001011" when "11011", -- t[27] = 11
         "0001010" when "11100", -- t[28] = 10
         "0001010" when "11101", -- t[29] = 10
         "0001001" when "11110", -- t[30] = 9
         "0001001" when "11111", -- t[31] = 9
         "-------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_2.
-- Decomposition:
--   alpha_2,2 = 2; sigma'_2,2 = 3; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t2_t2 is
  port ( a : in  std_logic_vector(1 downto 0);
         s : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of fp_log_log_18_t2_t2 is
  signal x : std_logic_vector(4 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0" when "00000", -- t[0] = 0
         "0" when "00001", -- t[1] = 0
         "0" when "00010", -- t[2] = 0
         "0" when "00011", -- t[3] = 0
         "0" when "00100", -- t[4] = 0
         "0" when "00101", -- t[5] = 0
         "0" when "00110", -- t[6] = 0
         "0" when "00111", -- t[7] = 0
         "0" when "01000", -- t[8] = 0
         "0" when "01001", -- t[9] = 0
         "0" when "01010", -- t[10] = 0
         "0" when "01011", -- t[11] = 0
         "0" when "01100", -- t[12] = 0
         "0" when "01101", -- t[13] = 0
         "0" when "01110", -- t[14] = 0
         "0" when "01111", -- t[15] = 0
         "0" when "10000", -- t[16] = 0
         "0" when "10001", -- t[17] = 0
         "0" when "10010", -- t[18] = 0
         "0" when "10011", -- t[19] = 0
         "0" when "10100", -- t[20] = 0
         "0" when "10101", -- t[21] = 0
         "0" when "10110", -- t[22] = 0
         "0" when "10111", -- t[23] = 0
         "0" when "11000", -- t[24] = 0
         "0" when "11001", -- t[25] = 0
         "0" when "11010", -- t[26] = 0
         "0" when "11011", -- t[27] = 0
         "0" when "11100", -- t[28] = 0
         "0" when "11101", -- t[29] = 0
         "0" when "11110", -- t[30] = 0
         "0" when "11111", -- t[31] = 0
         "-" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 5; beta_2 = 6; lambda_2 = 10;  m_2 = 2;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 5; rho_2,1 = 0; sigma_2,1 = 6; wO_2,1 = 7;
--   Q_2,2 (ROM):  alpha_2,2 = 2; rho_2,2 = 6; sigma_2,2 = 4; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_t2 is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(21 downto 0) );
end entity;

architecture arch of fp_log_log_18_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(4 downto 0);
  signal s      : std_logic_vector(9 downto 0);
  component fp_log_log_18_t2_pow is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  signal a_1    : std_logic_vector(4 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(4 downto 0);
  signal k_1    : std_logic_vector(6 downto 0);
  signal r0_1   : std_logic_vector(13 downto 0);
  signal r_1    : std_logic_vector(21 downto 0);
  component fp_log_log_18_t2_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  signal a_2    : std_logic_vector(1 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(2 downto 0);
  signal r0_2   : std_logic_vector(0 downto 0);
  signal r_2    : std_logic_vector(21 downto 0);
  component fp_log_log_18_t2_t2 is
    port ( a : in  std_logic_vector(1 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;
begin
  sign <= not b(5);
  b0 <= b(4 downto 0) xor (4 downto 0 => sign);

  pow : fp_log_log_18_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(4 downto 0);
  sign_1 <= not s(9);
  s_1 <= s(8 downto 4) xor (8 downto 4 => sign_1);
  t_1 : fp_log_log_18_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(6 downto 0) <=
    r0_1(13 downto 7) xor (13 downto 7 => ((sign_1)));
  r_1(21 downto 7) <= (21 downto 7 => ((sign_1)));

  a_2 <= a(4 downto 3);
  sign_2 <= not s(3);
  s_2 <= s(2 downto 0) xor (2 downto 0 => sign_2);
  t_2 : fp_log_log_18_t2_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(0 downto 0) <=
    r0_2 xor (0 downto 0 => ((sign_2)));
  r_2(21 downto 1) <= (21 downto 1 => ((sign_2)));

  r <= r_1 + r_2;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_fp_log.all;

entity fp_log_log_18_t2_clk is
  port ( a   : in  std_logic_vector(4 downto 0);
         b   : in  std_logic_vector(5 downto 0);
         r   : out std_logic_vector(21 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_18_t2_clk is
  signal sign_0 : std_logic;
  signal b0_0   : std_logic_vector(4 downto 0);
  signal s_0    : std_logic_vector(9 downto 0);
  component fp_log_log_18_t2_pow is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  signal a_1_0    : std_logic_vector(4 downto 0);
  signal sign_1_0 : std_logic;
  signal sign_1_1 : std_logic;
  signal sign_1_2 : std_logic;
  signal sign_1_3 : std_logic;
  signal s_1_0    : std_logic_vector(5 downto 0);
  signal s_1_1    : std_logic_vector(5 downto 0);
  signal k_1_0    : std_logic_vector(6 downto 0);
  signal k_1_1    : std_logic_vector(6 downto 0);
  signal r0_1_2   : std_logic_vector(12 downto 0);
  signal r1_1_2   : std_logic_vector(13 downto 0);
  signal r1_1_3   : std_logic_vector(13 downto 0);
  signal r_1_3    : std_logic_vector(21 downto 0);
  component fp_log_log_18_t2_t1 is
    port ( a : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  signal a_2_0    : std_logic_vector(1 downto 0);
  signal a_2_1    : std_logic_vector(1 downto 0);
  signal a_2_2    : std_logic_vector(1 downto 0);
  signal a_2_3    : std_logic_vector(1 downto 0);
  signal sign_2_0 : std_logic;
  signal sign_2_1 : std_logic;
  signal sign_2_2 : std_logic;
  signal sign_2_3 : std_logic;
  signal s_2_0    : std_logic_vector(2 downto 0);
  signal s_2_1    : std_logic_vector(2 downto 0);
  signal s_2_2    : std_logic_vector(2 downto 0);
  signal s_2_3    : std_logic_vector(2 downto 0);
  signal r0_2_3   : std_logic_vector(0 downto 0);
  signal r_2_3    : std_logic_vector(21 downto 0);
  component fp_log_log_18_t2_t2 is
    port ( a : in  std_logic_vector(1 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;
begin
  sign_0 <= not b(5);
  b0_0 <= b(4 downto 0) xor (4 downto 0 => sign_0);

  pow : fp_log_log_18_t2_pow
    port map ( x => b0_0,
               r => s_0 );

  a_1_0 <= a(4 downto 0);
  sign_1_0 <= not s_0(9);
  s_1_0 <= (s_0(8 downto 4) xor (8 downto 4 => sign_1_0)) & "1";
  t_1 : fp_log_log_18_t2_t1
    port map ( a => a_1_0,
               r => k_1_0 );

  mult_r0_1 : mult_clk
    generic map ( wX    => 7,
                  wY    => 6,
                  first => 0,
                  steps => 2 )
    port map ( nX  => k_1_1,
               nY  => s_1_1,
               nR  => r0_1_2,
               clk => clk );
  
  r1_1_2 <= "0" & r0_1_2;
  r_1_3(6 downto 0) <=
    r1_1_3(13 downto 7) xor (13 downto 7 => ((sign_1_3)));
  r_1_3(21 downto 7) <= (21 downto 7 => ((sign_1_3)));

  a_2_0 <= a(4 downto 3);
  sign_2_0 <= not s_0(3);
  s_2_0 <= s_0(2 downto 0) xor (2 downto 0 => sign_2_0);
  t_2 : fp_log_log_18_t2_t2
    port map ( a => a_2_3,
               s => s_2_3,
               r => r0_2_3 );
  r_2_3(0 downto 0) <=
    r0_2_3 xor (0 downto 0 => ((sign_2_3)));
  r_2_3(21 downto 1) <= (21 downto 1 => ((sign_2_3)));

  process(clk)
  begin
    if clk'event and clk = '1' then
      sign_1_1 <= sign_1_0;
      sign_1_2 <= sign_1_1;
      sign_1_3 <= sign_1_2;
      s_1_1    <= s_1_0;
      k_1_1    <= k_1_0;
      r1_1_3   <= r1_1_2;

      a_2_1    <= a_2_0;
      a_2_2    <= a_2_1;
      a_2_3    <= a_2_2;
      sign_2_1 <= sign_2_0;
      sign_2_2 <= sign_2_1;
      sign_2_3 <= sign_2_2;
      s_2_1    <= s_2_0;
      s_2_2    <= s_2_1;
      s_2_3    <= s_2_2;
    end if;
  end process;
  
  r <= r_1_3 + r_2_3;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18 is
  port ( x : in  std_logic_vector(17 downto 0);
         r : out std_logic_vector(21 downto 0) );
end entity;

architecture arch of fp_log_log_18 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(21 downto 0);
  component fp_log_log_18_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(21 downto 0) );
  end component;

  signal a_1 : std_logic_vector(6 downto 0);
  signal b_1 : std_logic_vector(10 downto 0);
  signal r_1 : std_logic_vector(21 downto 0);
  component fp_log_log_18_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(21 downto 0) );
  end component;

  signal a_2 : std_logic_vector(4 downto 0);
  signal b_2 : std_logic_vector(5 downto 0);
  signal r_2 : std_logic_vector(21 downto 0);
  component fp_log_log_18_t2 is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(21 downto 0) );
  end component;

begin
  a_0 <= x(17 downto 11);
  t_0 : fp_log_log_18_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(17 downto 11);
  b_1 <= x(10 downto 0);
  t_1 : fp_log_log_18_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(17 downto 13);
  b_2 <= x(10 downto 5);
  t_2 : fp_log_log_18_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_18_clk is
  port ( x   : in  std_logic_vector(17 downto 0);
         r   : out std_logic_vector(21 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_18_clk is
  signal x_0 : std_logic_vector(17 downto 0);
  signal x_1 : std_logic_vector(17 downto 0);
  signal x_2 : std_logic_vector(17 downto 0);
  signal x_3 : std_logic_vector(17 downto 0);
  
  signal a_0_3 : std_logic_vector(6 downto 0);
  signal r_0_3 : std_logic_vector(21 downto 0);
  signal r_0_4 : std_logic_vector(21 downto 0);
  component fp_log_log_18_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(21 downto 0) );
  end component;

  signal a_1_0 : std_logic_vector(6 downto 0);
  signal b_1_0 : std_logic_vector(10 downto 0);
  signal r_1_3 : std_logic_vector(21 downto 0);
  signal r_1_4 : std_logic_vector(21 downto 0);
  component fp_log_log_18_t1_clk is
    port ( a   : in  std_logic_vector(6 downto 0);
           b   : in  std_logic_vector(10 downto 0);
           r   : out std_logic_vector(21 downto 0);
           clk : in  std_logic );
  end component;

  signal a_2_0 : std_logic_vector(4 downto 0);
  signal b_2_0 : std_logic_vector(5 downto 0);
  signal r_2_3 : std_logic_vector(21 downto 0);
  signal r_2_4 : std_logic_vector(21 downto 0);
  component fp_log_log_18_t2_clk is
    port ( a   : in  std_logic_vector(4 downto 0);
           b   : in  std_logic_vector(5 downto 0);
           r   : out std_logic_vector(21 downto 0);
           clk : in  std_logic );
  end component;

begin
  x_0 <= x;
  
  a_0_3 <= x_3(17 downto 11);
  t_0 : fp_log_log_18_t0
    port map ( a => a_0_3,
               r => r_0_3 );

  a_1_0 <= x_0(17 downto 11);
  b_1_0 <= x_0(10 downto 0);
  t_1 : fp_log_log_18_t1_clk
    port map ( a   => a_1_0,
               b   => b_1_0,
               r   => r_1_3,
               clk => clk );

  a_2_0 <= x_0(17 downto 13);
  b_2_0 <= x_0(10 downto 5);
  t_2 : fp_log_log_18_t2_clk
    port map ( a   => a_2_0,
               b   => b_2_0,
               r         => r_2_3,
               clk => clk );

  process(clk)
  begin
    if clk'event and clk = '1' then
      x_1 <= x_0;
      x_2 <= x_1;
      x_3 <= x_2;
      r_0_4 <= r_0_3;
      r_1_4 <= r_1_3;
      r_2_4 <= r_2_3;
    end if;
  end process;
  
  r <= r_0_4 + r_1_4 + r_2_4;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 19; wO = 19.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 7; beta = 12;
--   T_0 (ROM):     alpha_0 = 7; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 7; beta_1 = 12;
--   T_2 (PowMult): alpha_2 = 6; beta_2 = 7.
-- Guard bits: g = 3.
-- Command line: logfp 19 19 2   rom 7 0   pm 7 12  ah 12 12 12  1 0  7 12 0   pm 6 7  ah 7 14 8  1 0  6 8 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 7; beta_0 = 0; wO_0 = 23.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19_t0 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(22 downto 0) );
end entity;

architecture arch of fp_log_log_19_t0 is
  signal x0   : std_logic_vector(6 downto 0);
  signal r0   : std_logic_vector(22 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110000110101011101000" when "0000000", -- t[0] = 5794536
          "10101111101000011010010" when "0000001", -- t[1] = 5755090
          "10101110011100110110010" when "0000010", -- t[2] = 5716402
          "10101101010010101100100" when "0000011", -- t[3] = 5678436
          "10101100001001111011100" when "0000100", -- t[4] = 5641180
          "10101011000010011111010" when "0000101", -- t[5] = 5604602
          "10101001111100010110001" when "0000110", -- t[6] = 5568689
          "10101000110111011100100" when "0000111", -- t[7] = 5533412
          "10100111110011110001001" when "0001000", -- t[8] = 5498761
          "10100110110001010000100" when "0001001", -- t[9] = 5464708
          "10100101101111111001100" when "0001010", -- t[10] = 5431244
          "10100100101111101001000" when "0001011", -- t[11] = 5398344
          "10100011110000011101111" when "0001100", -- t[12] = 5365999
          "10100010110010010101011" when "0001101", -- t[13] = 5334187
          "10100001110101001110010" when "0001110", -- t[14] = 5302898
          "10100000111001000110000" when "0001111", -- t[15] = 5272112
          "10011111111101111011110" when "0010000", -- t[16] = 5241822
          "10011111000011101100111" when "0010001", -- t[17] = 5212007
          "10011110001010011000110" when "0010010", -- t[18] = 5182662
          "10011101010001111100111" when "0010011", -- t[19] = 5153767
          "10011100011010011000101" when "0010100", -- t[20] = 5125317
          "10011011100011101001111" when "0010101", -- t[21] = 5097295
          "10011010101101101111110" when "0010110", -- t[22] = 5069694
          "10011001111000101000100" when "0010111", -- t[23] = 5042500
          "10011001000100010011011" when "0011000", -- t[24] = 5015707
          "10011000010000101110100" when "0011001", -- t[25] = 4989300
          "10010111011101111001011" when "0011010", -- t[26] = 4963275
          "10010110101011110010001" when "0011011", -- t[27] = 4937617
          "10010101111010011000010" when "0011100", -- t[28] = 4912322
          "10010101001001101010010" when "0011101", -- t[29] = 4887378
          "10010100011001100111100" when "0011110", -- t[30] = 4862780
          "10010011101010001110100" when "0011111", -- t[31] = 4838516
          "10010010111011011110110" when "0100000", -- t[32] = 4814582
          "10010010001101010110111" when "0100001", -- t[33] = 4790967
          "10010001011111110110100" when "0100010", -- t[34] = 4767668
          "10010000110010111100001" when "0100011", -- t[35] = 4744673
          "10010000000110100111100" when "0100100", -- t[36] = 4721980
          "10001111011010110111010" when "0100101", -- t[37] = 4699578
          "10001110101111101011001" when "0100110", -- t[38] = 4677465
          "10001110000101000001111" when "0100111", -- t[39] = 4655631
          "10001101011010111011000" when "0101000", -- t[40] = 4634072
          "10001100110001010101110" when "0101001", -- t[41] = 4612782
          "10001100001000010001011" when "0101010", -- t[42] = 4591755
          "10001011011111101101001" when "0101011", -- t[43] = 4570985
          "10001010110111101000101" when "0101100", -- t[44] = 4550469
          "10001010010000000010111" when "0101101", -- t[45] = 4530199
          "10001001101000111011100" when "0101110", -- t[46] = 4510172
          "10001001000010010001101" when "0101111", -- t[47] = 4490381
          "10001000011100000101000" when "0110000", -- t[48] = 4470824
          "10000111110110010100101" when "0110001", -- t[49] = 4451493
          "10000111010001000000100" when "0110010", -- t[50] = 4432388
          "10000110101100000111100" when "0110011", -- t[51] = 4413500
          "10000110000111101001100" when "0110100", -- t[52] = 4394828
          "10000101100011100101111" when "0110101", -- t[53] = 4376367
          "10000100111111111100001" when "0110110", -- t[54] = 4358113
          "10000100011100101011101" when "0110111", -- t[55] = 4340061
          "10000011111001110100001" when "0111000", -- t[56] = 4322209
          "10000011010111010100111" when "0111001", -- t[57] = 4304551
          "10000010110101001101111" when "0111010", -- t[58] = 4287087
          "10000010010011011110010" when "0111011", -- t[59] = 4269810
          "10000001110010000101111" when "0111100", -- t[60] = 4252719
          "10000001010001000100000" when "0111101", -- t[61] = 4235808
          "10000000110000011000101" when "0111110", -- t[62] = 4219077
          "10000000010000000011000" when "0111111", -- t[63] = 4202520
          "01111111110000000011000" when "1000000", -- t[64] = 4186136
          "01111111010000011000001" when "1000001", -- t[65] = 4169921
          "01111110110001000010001" when "1000010", -- t[66] = 4153873
          "01111110010010000000011" when "1000011", -- t[67] = 4137987
          "01111101110011010010111" when "1000100", -- t[68] = 4122263
          "01111101010100111001000" when "1000101", -- t[69] = 4106696
          "01111100110110110010100" when "1000110", -- t[70] = 4091284
          "01111100011000111111001" when "1000111", -- t[71] = 4076025
          "01111011111011011110101" when "1001000", -- t[72] = 4060917
          "01111011011110010000011" when "1001001", -- t[73] = 4045955
          "01111011000001010100100" when "1001010", -- t[74] = 4031140
          "01111010100100101010010" when "1001011", -- t[75] = 4016466
          "01111010001000010001110" when "1001100", -- t[76] = 4001934
          "01111001101100001010100" when "1001101", -- t[77] = 3987540
          "01111001010000010100010" when "1001110", -- t[78] = 3973282
          "01111000110100101110110" when "1001111", -- t[79] = 3959158
          "01111000011001011001110" when "1010000", -- t[80] = 3945166
          "01110111111110010100111" when "1010001", -- t[81] = 3931303
          "01110111100011100000001" when "1010010", -- t[82] = 3917569
          "01110111001000111011000" when "1010011", -- t[83] = 3903960
          "01110110101110100101100" when "1010100", -- t[84] = 3890476
          "01110110010100011111001" when "1010101", -- t[85] = 3877113
          "01110101111010100111110" when "1010110", -- t[86] = 3863870
          "01110101100000111111010" when "1010111", -- t[87] = 3850746
          "01110101000111100101011" when "1011000", -- t[88] = 3837739
          "01110100101110011001110" when "1011001", -- t[89] = 3824846
          "01110100010101011100010" when "1011010", -- t[90] = 3812066
          "01110011111100101100110" when "1011011", -- t[91] = 3799398
          "01110011100100001011000" when "1011100", -- t[92] = 3786840
          "01110011001011110110110" when "1011101", -- t[93] = 3774390
          "01110010110011110000000" when "1011110", -- t[94] = 3762048
          "01110010011011110110010" when "1011111", -- t[95] = 3749810
          "01110010000100001001100" when "1100000", -- t[96] = 3737676
          "01110001101100101001100" when "1100001", -- t[97] = 3725644
          "01110001010101010110010" when "1100010", -- t[98] = 3713714
          "01110000111110001111010" when "1100011", -- t[99] = 3701882
          "01110000100111010100101" when "1100100", -- t[100] = 3690149
          "01110000010000100110000" when "1100101", -- t[101] = 3678512
          "01101111111010000011011" when "1100110", -- t[102] = 3666971
          "01101111100011101100100" when "1100111", -- t[103] = 3655524
          "01101111001101100001001" when "1101000", -- t[104] = 3644169
          "01101110110111100001010" when "1101001", -- t[105] = 3632906
          "01101110100001101100110" when "1101010", -- t[106] = 3621734
          "01101110001100000011010" when "1101011", -- t[107] = 3610650
          "01101101110110100100111" when "1101100", -- t[108] = 3599655
          "01101101100001010001010" when "1101101", -- t[109] = 3588746
          "01101101001100001000011" when "1101110", -- t[110] = 3577923
          "01101100110111001010001" when "1101111", -- t[111] = 3567185
          "01101100100010010110010" when "1110000", -- t[112] = 3556530
          "01101100001101101100101" when "1110001", -- t[113] = 3545957
          "01101011111001001101010" when "1110010", -- t[114] = 3535466
          "01101011100100110111110" when "1110011", -- t[115] = 3525054
          "01101011010000101100010" when "1110100", -- t[116] = 3514722
          "01101010111100101010101" when "1110101", -- t[117] = 3504469
          "01101010101000110010100" when "1110110", -- t[118] = 3494292
          "01101010010101000100000" when "1110111", -- t[119] = 3484192
          "01101010000001011110111" when "1111000", -- t[120] = 3474167
          "01101001101110000011001" when "1111001", -- t[121] = 3464217
          "01101001011010110000100" when "1111010", -- t[122] = 3454340
          "01101001000111100110111" when "1111011", -- t[123] = 3444535
          "01101000110100100110010" when "1111100", -- t[124] = 3434802
          "01101000100001101110100" when "1111101", -- t[125] = 3425140
          "01101000001110111111101" when "1111110", -- t[126] = 3415549
          "01100111111100011001010" when "1111111", -- t[127] = 3406026
          "-----------------------" when others;

  r(22 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 12; mu_1 = 12; lambda_1 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19_t1_pow is
  port ( x : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_19_t1_pow is
  signal pp0 : std_logic_vector(10 downto 0);
  signal r0 : std_logic_vector(10 downto 0);
begin
  pp0(10) <= x(10);

  pp0(9) <= x(9);

  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(10 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 7; wO_1,1 = 16.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19_t1_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of fp_log_log_19_t1_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "1001101110010100" when "0000000", -- t[0] = 39828
         "1001100010011000" when "0000001", -- t[1] = 39064
         "1001010110110100" when "0000010", -- t[2] = 38324
         "1001001011101000" when "0000011", -- t[3] = 37608
         "1001000000110010" when "0000100", -- t[4] = 36914
         "1000110110010011" when "0000101", -- t[5] = 36243
         "1000101100001000" when "0000110", -- t[6] = 35592
         "1000100010010001" when "0000111", -- t[7] = 34961
         "1000011000101101" when "0001000", -- t[8] = 34349
         "1000001111011100" when "0001001", -- t[9] = 33756
         "1000000110011100" when "0001010", -- t[10] = 33180
         "0111111101101100" when "0001011", -- t[11] = 32620
         "0111110101001101" when "0001100", -- t[12] = 32077
         "0111101100111101" when "0001101", -- t[13] = 31549
         "0111100100111011" when "0001110", -- t[14] = 31035
         "0111011101001000" when "0001111", -- t[15] = 30536
         "0111010101100011" when "0010000", -- t[16] = 30051
         "0111001110001010" when "0010001", -- t[17] = 29578
         "0111000110111110" when "0010010", -- t[18] = 29118
         "0110111111111111" when "0010011", -- t[19] = 28671
         "0110111001001011" when "0010100", -- t[20] = 28235
         "0110110010100010" when "0010101", -- t[21] = 27810
         "0110101100000100" when "0010110", -- t[22] = 27396
         "0110100101110000" when "0010111", -- t[23] = 26992
         "0110011111100111" when "0011000", -- t[24] = 26599
         "0110011001100111" when "0011001", -- t[25] = 26215
         "0110010011110000" when "0011010", -- t[26] = 25840
         "0110001110000011" when "0011011", -- t[27] = 25475
         "0110001000011110" when "0011100", -- t[28] = 25118
         "0110000011000010" when "0011101", -- t[29] = 24770
         "0101111101101110" when "0011110", -- t[30] = 24430
         "0101111000100010" when "0011111", -- t[31] = 24098
         "0101110011011101" when "0100000", -- t[32] = 23773
         "0101101110100000" when "0100001", -- t[33] = 23456
         "0101101001101010" when "0100010", -- t[34] = 23146
         "0101100100111011" when "0100011", -- t[35] = 22843
         "0101100000010011" when "0100100", -- t[36] = 22547
         "0101011011110001" when "0100101", -- t[37] = 22257
         "0101010111010101" when "0100110", -- t[38] = 21973
         "0101010010111111" when "0100111", -- t[39] = 21695
         "0101001110110000" when "0101000", -- t[40] = 21424
         "0101001010100110" when "0101001", -- t[41] = 21158
         "0101000110100001" when "0101010", -- t[42] = 20897
         "0101000010100010" when "0101011", -- t[43] = 20642
         "0100111110101001" when "0101100", -- t[44] = 20393
         "0100111010110100" when "0101101", -- t[45] = 20148
         "0100110111000100" when "0101110", -- t[46] = 19908
         "0100110011011001" when "0101111", -- t[47] = 19673
         "0100101111110011" when "0110000", -- t[48] = 19443
         "0100101100010001" when "0110001", -- t[49] = 19217
         "0100101000110100" when "0110010", -- t[50] = 18996
         "0100100101011011" when "0110011", -- t[51] = 18779
         "0100100010000110" when "0110100", -- t[52] = 18566
         "0100011110110101" when "0110101", -- t[53] = 18357
         "0100011011101000" when "0110110", -- t[54] = 18152
         "0100011000011111" when "0110111", -- t[55] = 17951
         "0100010101011010" when "0111000", -- t[56] = 17754
         "0100010010011000" when "0111001", -- t[57] = 17560
         "0100001111011010" when "0111010", -- t[58] = 17370
         "0100001100100000" when "0111011", -- t[59] = 17184
         "0100001001101000" when "0111100", -- t[60] = 17000
         "0100000110110100" when "0111101", -- t[61] = 16820
         "0100000100000100" when "0111110", -- t[62] = 16644
         "0100000001010110" when "0111111", -- t[63] = 16470
         "0011111110101011" when "1000000", -- t[64] = 16299
         "0011111100000011" when "1000001", -- t[65] = 16131
         "0011111001011111" when "1000010", -- t[66] = 15967
         "0011110110111101" when "1000011", -- t[67] = 15805
         "0011110100011101" when "1000100", -- t[68] = 15645
         "0011110010000001" when "1000101", -- t[69] = 15489
         "0011101111100111" when "1000110", -- t[70] = 15335
         "0011101101010000" when "1000111", -- t[71] = 15184
         "0011101010111011" when "1001000", -- t[72] = 15035
         "0011101000101000" when "1001001", -- t[73] = 14888
         "0011100110011000" when "1001010", -- t[74] = 14744
         "0011100100001010" when "1001011", -- t[75] = 14602
         "0011100001111111" when "1001100", -- t[76] = 14463
         "0011011111110110" when "1001101", -- t[77] = 14326
         "0011011101101111" when "1001110", -- t[78] = 14191
         "0011011011101010" when "1001111", -- t[79] = 14058
         "0011011001100111" when "1010000", -- t[80] = 13927
         "0011010111100110" when "1010001", -- t[81] = 13798
         "0011010101100111" when "1010010", -- t[82] = 13671
         "0011010011101010" when "1010011", -- t[83] = 13546
         "0011010001110000" when "1010100", -- t[84] = 13424
         "0011001111110110" when "1010101", -- t[85] = 13302
         "0011001101111111" when "1010110", -- t[86] = 13183
         "0011001100001010" when "1010111", -- t[87] = 13066
         "0011001010010110" when "1011000", -- t[88] = 12950
         "0011001000100100" when "1011001", -- t[89] = 12836
         "0011000110110100" when "1011010", -- t[90] = 12724
         "0011000101000101" when "1011011", -- t[91] = 12613
         "0011000011011000" when "1011100", -- t[92] = 12504
         "0011000001101100" when "1011101", -- t[93] = 12396
         "0011000000000010" when "1011110", -- t[94] = 12290
         "0010111110011010" when "1011111", -- t[95] = 12186
         "0010111100110011" when "1100000", -- t[96] = 12083
         "0010111011001101" when "1100001", -- t[97] = 11981
         "0010111001101001" when "1100010", -- t[98] = 11881
         "0010111000000110" when "1100011", -- t[99] = 11782
         "0010110110100101" when "1100100", -- t[100] = 11685
         "0010110101000101" when "1100101", -- t[101] = 11589
         "0010110011100110" when "1100110", -- t[102] = 11494
         "0010110010001001" when "1100111", -- t[103] = 11401
         "0010110000101100" when "1101000", -- t[104] = 11308
         "0010101111010001" when "1101001", -- t[105] = 11217
         "0010101101111000" when "1101010", -- t[106] = 11128
         "0010101100011111" when "1101011", -- t[107] = 11039
         "0010101011001000" when "1101100", -- t[108] = 10952
         "0010101001110010" when "1101101", -- t[109] = 10866
         "0010101000011101" when "1101110", -- t[110] = 10781
         "0010100111001001" when "1101111", -- t[111] = 10697
         "0010100101110110" when "1110000", -- t[112] = 10614
         "0010100100100100" when "1110001", -- t[113] = 10532
         "0010100011010011" when "1110010", -- t[114] = 10451
         "0010100010000011" when "1110011", -- t[115] = 10371
         "0010100000110101" when "1110100", -- t[116] = 10293
         "0010011111100111" when "1110101", -- t[117] = 10215
         "0010011110011010" when "1110110", -- t[118] = 10138
         "0010011101001110" when "1110111", -- t[119] = 10062
         "0010011100000100" when "1111000", -- t[120] = 9988
         "0010011010111010" when "1111001", -- t[121] = 9914
         "0010011001110001" when "1111010", -- t[122] = 9841
         "0010011000101000" when "1111011", -- t[123] = 9768
         "0010010111100001" when "1111100", -- t[124] = 9697
         "0010010110011011" when "1111101", -- t[125] = 9627
         "0010010101010101" when "1111110", -- t[126] = 9557
         "0010010100010001" when "1111111", -- t[127] = 9489
         "----------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 7; beta_1 = 12; lambda_1 = 12;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 7; rho_1,1 = 0; sigma_1,1 = 12; wO_1,1 = 16.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(22 downto 0) );
end entity;

architecture arch of fp_log_log_19_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(10 downto 0);
  signal s      : std_logic_vector(11 downto 0);
  component fp_log_log_19_t1_pow is
    port ( x : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(10 downto 0);
  signal k_1    : std_logic_vector(15 downto 0);
  signal r0_1   : std_logic_vector(28 downto 0);
  signal r_1    : std_logic_vector(22 downto 0);
  component fp_log_log_19_t1_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(15 downto 0) );
  end component;
begin
  sign <= not b(11);
  b0 <= b(10 downto 0) xor (10 downto 0 => sign);

  pow : fp_log_log_19_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(11);
  s_1 <= s(10 downto 0) xor (10 downto 0 => sign_1);
  t_1 : fp_log_log_19_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(15 downto 0) <=
    r0_1(28 downto 13) xor (28 downto 13 => (not (sign xor sign_1)));
  r_1(22 downto 16) <= (22 downto 16 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 7; mu_2 = 14; lambda_2 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19_t2_pow is
  port ( x : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_log_log_19_t2_pow is
  signal pp0 : std_logic_vector(12 downto 0);
  signal pp1 : std_logic_vector(12 downto 0);
  signal pp2 : std_logic_vector(12 downto 0);
  signal pp3 : std_logic_vector(12 downto 0);
  signal r0 : std_logic_vector(12 downto 0);
begin
  pp0(12) <= '0';
  pp1(12) <= '0';
  pp2(12) <= '0';
  pp3(12) <= '0';

  pp0(11) <= x(4) and x(5);
  pp1(11) <= x(5);
  pp2(11) <= '0';
  pp3(11) <= '0';

  pp0(10) <= x(3) and x(5);
  pp1(10) <= '0';
  pp2(10) <= '0';
  pp3(10) <= '0';

  pp0(9) <= x(2) and x(5);
  pp1(9) <= x(3) and x(4);
  pp2(9) <= x(4);
  pp3(9) <= '0';

  pp0(8) <= x(1) and x(5);
  pp1(8) <= x(2) and x(4);
  pp2(8) <= '0';
  pp3(8) <= '0';

  pp0(7) <= x(0) and x(5);
  pp1(7) <= x(1) and x(4);
  pp2(7) <= x(2) and x(3);
  pp3(7) <= x(3);

  pp0(6) <= x(0) and x(4);
  pp1(6) <= x(1) and x(3);
  pp2(6) <= x(5);
  pp3(6) <= '0';

  pp0(5) <= x(0) and x(3);
  pp1(5) <= x(1) and x(2);
  pp2(5) <= x(2);
  pp3(5) <= x(4);

  pp0(4) <= x(0) and x(2);
  pp1(4) <= x(3);
  pp2(4) <= '0';
  pp3(4) <= '0';

  pp0(3) <= x(0) and x(1);
  pp1(3) <= x(1);
  pp2(3) <= x(2);
  pp3(3) <= '0';

  pp0(2) <= x(0);
  pp1(2) <= x(1);
  pp2(2) <= '0';
  pp3(2) <= '0';

  pp0(1) <= '0';
  pp1(1) <= '0';
  pp2(1) <= '0';
  pp3(1) <= '0';

  pp0(0) <= '0';
  pp1(0) <= '0';
  pp2(0) <= '0';
  pp3(0) <= '0';

  r0 <= pp0 + pp1 + pp2 + pp3;
  r <= "1" & r0(12 downto 6);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 6; wO_2,1 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19_t2_t1 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_log_log_19_t2_t1 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a;

  with x select
    r <= "10111111" when "000000", -- t[0] = 191
         "10110011" when "000001", -- t[1] = 179
         "10101000" when "000010", -- t[2] = 168
         "10011110" when "000011", -- t[3] = 158
         "10010100" when "000100", -- t[4] = 148
         "10001100" when "000101", -- t[5] = 140
         "10000100" when "000110", -- t[6] = 132
         "01111101" when "000111", -- t[7] = 125
         "01110110" when "001000", -- t[8] = 118
         "01110000" when "001001", -- t[9] = 112
         "01101010" when "001010", -- t[10] = 106
         "01100101" when "001011", -- t[11] = 101
         "01100000" when "001100", -- t[12] = 96
         "01011011" when "001101", -- t[13] = 91
         "01010111" when "001110", -- t[14] = 87
         "01010011" when "001111", -- t[15] = 83
         "01001111" when "010000", -- t[16] = 79
         "01001100" when "010001", -- t[17] = 76
         "01001000" when "010010", -- t[18] = 72
         "01000101" when "010011", -- t[19] = 69
         "01000010" when "010100", -- t[20] = 66
         "01000000" when "010101", -- t[21] = 64
         "00111101" when "010110", -- t[22] = 61
         "00111011" when "010111", -- t[23] = 59
         "00111000" when "011000", -- t[24] = 56
         "00110110" when "011001", -- t[25] = 54
         "00110100" when "011010", -- t[26] = 52
         "00110010" when "011011", -- t[27] = 50
         "00110000" when "011100", -- t[28] = 48
         "00101111" when "011101", -- t[29] = 47
         "00101101" when "011110", -- t[30] = 45
         "00101011" when "011111", -- t[31] = 43
         "00101010" when "100000", -- t[32] = 42
         "00101001" when "100001", -- t[33] = 41
         "00100111" when "100010", -- t[34] = 39
         "00100110" when "100011", -- t[35] = 38
         "00100101" when "100100", -- t[36] = 37
         "00100011" when "100101", -- t[37] = 35
         "00100010" when "100110", -- t[38] = 34
         "00100001" when "100111", -- t[39] = 33
         "00100000" when "101000", -- t[40] = 32
         "00011111" when "101001", -- t[41] = 31
         "00011110" when "101010", -- t[42] = 30
         "00011101" when "101011", -- t[43] = 29
         "00011101" when "101100", -- t[44] = 29
         "00011100" when "101101", -- t[45] = 28
         "00011011" when "101110", -- t[46] = 27
         "00011010" when "101111", -- t[47] = 26
         "00011001" when "110000", -- t[48] = 25
         "00011001" when "110001", -- t[49] = 25
         "00011000" when "110010", -- t[50] = 24
         "00010111" when "110011", -- t[51] = 23
         "00010111" when "110100", -- t[52] = 23
         "00010110" when "110101", -- t[53] = 22
         "00010110" when "110110", -- t[54] = 22
         "00010101" when "110111", -- t[55] = 21
         "00010100" when "111000", -- t[56] = 20
         "00010100" when "111001", -- t[57] = 20
         "00010011" when "111010", -- t[58] = 19
         "00010011" when "111011", -- t[59] = 19
         "00010010" when "111100", -- t[60] = 18
         "00010010" when "111101", -- t[61] = 18
         "00010010" when "111110", -- t[62] = 18
         "00010001" when "111111", -- t[63] = 17
         "--------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 6; beta_2 = 7; lambda_2 = 8;  m_2 = 1;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 6; rho_2,1 = 0; sigma_2,1 = 8; wO_2,1 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19_t2 is
  port ( a : in  std_logic_vector(5 downto 0);
         b : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(22 downto 0) );
end entity;

architecture arch of fp_log_log_19_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(5 downto 0);
  signal s      : std_logic_vector(7 downto 0);
  component fp_log_log_19_t2_pow is
    port ( x : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  signal a_1    : std_logic_vector(5 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(6 downto 0);
  signal k_1    : std_logic_vector(7 downto 0);
  signal r0_1   : std_logic_vector(16 downto 0);
  signal r_1    : std_logic_vector(22 downto 0);
  component fp_log_log_19_t2_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;
begin
  sign <= not b(6);
  b0 <= b(5 downto 0) xor (5 downto 0 => sign);

  pow : fp_log_log_19_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(5 downto 0);
  sign_1 <= not s(7);
  s_1 <= s(6 downto 0) xor (6 downto 0 => sign_1);
  t_1 : fp_log_log_19_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(7 downto 0) <=
    r0_1(16 downto 9) xor (16 downto 9 => ((sign_1)));
  r_1(22 downto 8) <= (22 downto 8 => ((sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_19 is
  port ( x : in  std_logic_vector(18 downto 0);
         r : out std_logic_vector(22 downto 0) );
end entity;

architecture arch of fp_log_log_19 is
  signal a_0 : std_logic_vector(6 downto 0);
  signal r_0 : std_logic_vector(22 downto 0);
  component fp_log_log_19_t0 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(22 downto 0) );
  end component;

  signal a_1 : std_logic_vector(6 downto 0);
  signal b_1 : std_logic_vector(11 downto 0);
  signal r_1 : std_logic_vector(22 downto 0);
  component fp_log_log_19_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(22 downto 0) );
  end component;

  signal a_2 : std_logic_vector(5 downto 0);
  signal b_2 : std_logic_vector(6 downto 0);
  signal r_2 : std_logic_vector(22 downto 0);
  component fp_log_log_19_t2 is
    port ( a : in  std_logic_vector(5 downto 0);
           b : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(22 downto 0) );
  end component;

begin
  a_0 <= x(18 downto 12);
  t_0 : fp_log_log_19_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(18 downto 12);
  b_1 <= x(11 downto 0);
  t_1 : fp_log_log_19_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(18 downto 13);
  b_2 <= x(11 downto 5);
  t_2 : fp_log_log_19_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 20; wO = 20.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 8; beta = 12;
--   T_0 (ROM):     alpha_0 = 8; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 8; beta_1 = 12;
--   T_2 (PowMult): alpha_2 = 6; beta_2 = 6.
-- Guard bits: g = 3.
-- Command line: logfp 20 20 2   rom 8 0   pm 8 12  ah 12 12 12  1 0  8 12 0   pm 6 6  ah 6 12 8  1 0  6 8 0


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 8; beta_0 = 0; wO_0 = 24.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20_t0 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(23 downto 0) );
end entity;

architecture arch of fp_log_log_20_t0 is
  signal x0   : std_logic_vector(7 downto 0);
  signal r0   : std_logic_vector(23 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "101100010010001111000010" when "00000000", -- t[0] = 11609026
          "101100001000100000101110" when "00000001", -- t[1] = 11569198
          "101011111110111000011011" when "00000010", -- t[2] = 11529755
          "101011110101010110000011" when "00000011", -- t[3] = 11490691
          "101011101011111001100011" when "00000100", -- t[4] = 11452003
          "101011100010100010101111" when "00000101", -- t[5] = 11413679
          "101011011001010001100100" when "00000110", -- t[6] = 11375716
          "101011010000000101111101" when "00000111", -- t[7] = 11338109
          "101011000110111111110101" when "00001000", -- t[8] = 11300853
          "101010111101111111000011" when "00001001", -- t[9] = 11263939
          "101010110101000011100010" when "00001010", -- t[10] = 11227362
          "101010101100001101010000" when "00001011", -- t[11] = 11191120
          "101010100011011100000111" when "00001100", -- t[12] = 11155207
          "101010011010101111111111" when "00001101", -- t[13] = 11119615
          "101010010010001000110100" when "00001110", -- t[14] = 11084340
          "101010001001100110100011" when "00001111", -- t[15] = 11049379
          "101010000001001001001000" when "00010000", -- t[16] = 11014728
          "101001111000110000011010" when "00010001", -- t[17] = 10980378
          "101001110000011100010111" when "00010010", -- t[18] = 10946327
          "101001101000001100111011" when "00010011", -- t[19] = 10912571
          "101001100000000010000100" when "00010100", -- t[20] = 10879108
          "101001010111111011101000" when "00010101", -- t[21] = 10845928
          "101001001111111001100110" when "00010110", -- t[22] = 10813030
          "101001000111111011111010" when "00010111", -- t[23] = 10780410
          "101001000000000010100001" when "00011000", -- t[24] = 10748065
          "101000111000001101010100" when "00011001", -- t[25] = 10715988
          "101000110000011100010001" when "00011010", -- t[26] = 10684177
          "101000101000101111010100" when "00011011", -- t[27] = 10652628
          "101000100001000110011011" when "00011100", -- t[28] = 10621339
          "101000011001100001100000" when "00011101", -- t[29] = 10590304
          "101000010010000000100000" when "00011110", -- t[30] = 10559520
          "101000001010100011010111" when "00011111", -- t[31] = 10528983
          "101000000011001010000101" when "00100000", -- t[32] = 10498693
          "100111111011110100100010" when "00100001", -- t[33] = 10468642
          "100111110100100010101101" when "00100010", -- t[34] = 10438829
          "100111101101010100100011" when "00100011", -- t[35] = 10409251
          "100111100110001010000001" when "00100100", -- t[36] = 10379905
          "100111011111000011000011" when "00100101", -- t[37] = 10350787
          "100111010111111111100110" when "00100110", -- t[38] = 10321894
          "100111010000111111100111" when "00100111", -- t[39] = 10293223
          "100111001010000011000101" when "00101000", -- t[40] = 10264773
          "100111000011001001111010" when "00101001", -- t[41] = 10236538
          "100110111100010100000101" when "00101010", -- t[42] = 10208517
          "100110110101100001100011" when "00101011", -- t[43] = 10180707
          "100110101110110010010011" when "00101100", -- t[44] = 10153107
          "100110101000000110001111" when "00101101", -- t[45] = 10125711
          "100110100001011101010110" when "00101110", -- t[46] = 10098518
          "100110011010110111100110" when "00101111", -- t[47] = 10071526
          "100110010100010100111101" when "00110000", -- t[48] = 10044733
          "100110001101110101010110" when "00110001", -- t[49] = 10018134
          "100110000111011000110000" when "00110010", -- t[50] = 9991728
          "100110000000111111001010" when "00110011", -- t[51] = 9965514
          "100101111010101000100000" when "00110100", -- t[52] = 9939488
          "100101110100010100110000" when "00110101", -- t[53] = 9913648
          "100101101110000011110111" when "00110110", -- t[54] = 9887991
          "100101100111110101110100" when "00110111", -- t[55] = 9862516
          "100101100001101010100101" when "00111000", -- t[56] = 9837221
          "100101011011100010000111" when "00111001", -- t[57] = 9812103
          "100101010101011100010111" when "00111010", -- t[58] = 9787159
          "100101001111011001010101" when "00111011", -- t[59] = 9762389
          "100101001001011000111111" when "00111100", -- t[60] = 9737791
          "100101000011011011010001" when "00111101", -- t[61] = 9713361
          "100100111101100000001010" when "00111110", -- t[62] = 9689098
          "100100110111100111101000" when "00111111", -- t[63] = 9665000
          "100100110001110001101010" when "01000000", -- t[64] = 9641066
          "100100101011111110001100" when "01000001", -- t[65] = 9617292
          "100100100110001101001111" when "01000010", -- t[66] = 9593679
          "100100100000011110101110" when "01000011", -- t[67] = 9570222
          "100100011010110010101011" when "01000100", -- t[68] = 9546923
          "100100010101001001000001" when "01000101", -- t[69] = 9523777
          "100100001111100001101111" when "01000110", -- t[70] = 9500783
          "100100001001111100110100" when "01000111", -- t[71] = 9477940
          "100100000100011010001111" when "01001000", -- t[72] = 9455247
          "100011111110111001111100" when "01001001", -- t[73] = 9432700
          "100011111001011011111011" when "01001010", -- t[74] = 9410299
          "100011110100000000001011" when "01001011", -- t[75] = 9388043
          "100011101110100110101001" when "01001100", -- t[76] = 9365929
          "100011101001001111010100" when "01001101", -- t[77] = 9343956
          "100011100011111010001011" when "01001110", -- t[78] = 9322123
          "100011011110100111001100" when "01001111", -- t[79] = 9300428
          "100011011001010110010101" when "01010000", -- t[80] = 9278869
          "100011010100000111100110" when "01010001", -- t[81] = 9257446
          "100011001110111010111100" when "01010010", -- t[82] = 9236156
          "100011001001110000010110" when "01010011", -- t[83] = 9214998
          "100011000100100111110100" when "01010100", -- t[84] = 9193972
          "100010111111100001010010" when "01010101", -- t[85] = 9173074
          "100010111010011100110001" when "01010110", -- t[86] = 9152305
          "100010110101011010001110" when "01010111", -- t[87] = 9131662
          "100010110000011001101010" when "01011000", -- t[88] = 9111146
          "100010101011011011000001" when "01011001", -- t[89] = 9090753
          "100010100110011110010100" when "01011010", -- t[90] = 9070484
          "100010100001100011011111" when "01011011", -- t[91] = 9050335
          "100010011100101010100100" when "01011100", -- t[92] = 9030308
          "100010010111110011100000" when "01011101", -- t[93] = 9010400
          "100010010010111110010010" when "01011110", -- t[94] = 8990610
          "100010001110001010111000" when "01011111", -- t[95] = 8970936
          "100010001001011001010011" when "01100000", -- t[96] = 8951379
          "100010000100101001100000" when "01100001", -- t[97] = 8931936
          "100001111111111011011110" when "01100010", -- t[98] = 8912606
          "100001111011001111001101" when "01100011", -- t[99] = 8893389
          "100001110110100100101011" when "01100100", -- t[100] = 8874283
          "100001110001111011110111" when "01100101", -- t[101] = 8855287
          "100001101101010100110000" when "01100110", -- t[102] = 8836400
          "100001101000101111010101" when "01100111", -- t[103] = 8817621
          "100001100100001011100101" when "01101000", -- t[104] = 8798949
          "100001011111101001011111" when "01101001", -- t[105] = 8780383
          "100001011011001001000010" when "01101010", -- t[106] = 8761922
          "100001010110101010001101" when "01101011", -- t[107] = 8743565
          "100001010010001100111111" when "01101100", -- t[108] = 8725311
          "100001001101110001010110" when "01101101", -- t[109] = 8707158
          "100001001001010111010011" when "01101110", -- t[110] = 8689107
          "100001000100111110110011" when "01101111", -- t[111] = 8671155
          "100001000000100111110111" when "01110000", -- t[112] = 8653303
          "100000111100010010011101" when "01110001", -- t[113] = 8635549
          "100000110111111110100100" when "01110010", -- t[114] = 8617892
          "100000110011101100001100" when "01110011", -- t[115] = 8600332
          "100000101111011011010011" when "01110100", -- t[116] = 8582867
          "100000101011001011111001" when "01110101", -- t[117] = 8565497
          "100000100110111101111100" when "01110110", -- t[118] = 8548220
          "100000100010110001011100" when "01110111", -- t[119] = 8531036
          "100000011110100110011001" when "01111000", -- t[120] = 8513945
          "100000011010011100110001" when "01111001", -- t[121] = 8496945
          "100000010110010100100011" when "01111010", -- t[122] = 8480035
          "100000010010001101101110" when "01111011", -- t[123] = 8463214
          "100000001110001000010011" when "01111100", -- t[124] = 8446483
          "100000001010000100010000" when "01111101", -- t[125] = 8429840
          "100000000110000001100011" when "01111110", -- t[126] = 8413283
          "100000000010000000001110" when "01111111", -- t[127] = 8396814
          "011111111110000000001110" when "10000000", -- t[128] = 8380430
          "011111111010000001100011" when "10000001", -- t[129] = 8364131
          "011111110110000100001100" when "10000010", -- t[130] = 8347916
          "011111110010001000001000" when "10000011", -- t[131] = 8331784
          "011111101110001101011000" when "10000100", -- t[132] = 8315736
          "011111101010010011111001" when "10000101", -- t[133] = 8299769
          "011111100110011011101100" when "10000110", -- t[134] = 8283884
          "011111100010100100101111" when "10000111", -- t[135] = 8268079
          "011111011110101111000011" when "10001000", -- t[136] = 8252355
          "011111011010111010100110" when "10001001", -- t[137] = 8236710
          "011111010111000111010111" when "10001010", -- t[138] = 8221143
          "011111010011010101010110" when "10001011", -- t[139] = 8205654
          "011111001111100100100011" when "10001100", -- t[140] = 8190243
          "011111001011110100111100" when "10001101", -- t[141] = 8174908
          "011111001000000110100001" when "10001110", -- t[142] = 8159649
          "011111000100011001010001" when "10001111", -- t[143] = 8144465
          "011111000000101101001101" when "10010000", -- t[144] = 8129357
          "011110111101000010010010" when "10010001", -- t[145] = 8114322
          "011110111001011000100001" when "10010010", -- t[146] = 8099361
          "011110110101101111111001" when "10010011", -- t[147] = 8084473
          "011110110010001000011001" when "10010100", -- t[148] = 8069657
          "011110101110100010000001" when "10010101", -- t[149] = 8054913
          "011110101010111100110000" when "10010110", -- t[150] = 8040240
          "011110100111011000100110" when "10010111", -- t[151] = 8025638
          "011110100011110101100010" when "10011000", -- t[152] = 8011106
          "011110100000010011100011" when "10011001", -- t[153] = 7996643
          "011110011100110010101001" when "10011010", -- t[154] = 7982249
          "011110011001010010110011" when "10011011", -- t[155] = 7967923
          "011110010101110100000001" when "10011100", -- t[156] = 7953665
          "011110010010010110010010" when "10011101", -- t[157] = 7939474
          "011110001110111001100110" when "10011110", -- t[158] = 7925350
          "011110001011011101111101" when "10011111", -- t[159] = 7911293
          "011110001000000011010101" when "10100000", -- t[160] = 7897301
          "011110000100101001101110" when "10100001", -- t[161] = 7883374
          "011110000001010001000111" when "10100010", -- t[162] = 7869511
          "011101111101111001100001" when "10100011", -- t[163] = 7855713
          "011101111010100010111011" when "10100100", -- t[164] = 7841979
          "011101110111001101010100" when "10100101", -- t[165] = 7828308
          "011101110011111000101011" when "10100110", -- t[166] = 7814699
          "011101110000100101000000" when "10100111", -- t[167] = 7801152
          "011101101101010010010100" when "10101000", -- t[168] = 7787668
          "011101101010000000100100" when "10101001", -- t[169] = 7774244
          "011101100110101111110010" when "10101010", -- t[170] = 7760882
          "011101100011011111111011" when "10101011", -- t[171] = 7747579
          "011101100000010001000001" when "10101100", -- t[172] = 7734337
          "011101011101000011000010" when "10101101", -- t[173] = 7721154
          "011101011001110101111101" when "10101110", -- t[174] = 7708029
          "011101010110101001110100" when "10101111", -- t[175] = 7694964
          "011101010011011110100100" when "10110000", -- t[176] = 7681956
          "011101010000010100001111" when "10110001", -- t[177] = 7669007
          "011101001101001010110010" when "10110010", -- t[178] = 7656114
          "011101001010000010001110" when "10110011", -- t[179] = 7643278
          "011101000110111010100011" when "10110100", -- t[180] = 7630499
          "011101000011110011101111" when "10110101", -- t[181] = 7617775
          "011101000000101101110011" when "10110110", -- t[182] = 7605107
          "011100111101101000101110" when "10110111", -- t[183] = 7592494
          "011100111010100100100001" when "10111000", -- t[184] = 7579937
          "011100110111100001001001" when "10111001", -- t[185] = 7567433
          "011100110100011110100111" when "10111010", -- t[186] = 7554983
          "011100110001011100111011" when "10111011", -- t[187] = 7542587
          "011100101110011100000100" when "10111100", -- t[188] = 7530244
          "011100101011011100000010" when "10111101", -- t[189] = 7517954
          "011100101000011100110101" when "10111110", -- t[190] = 7505717
          "011100100101011110011011" when "10111111", -- t[191] = 7493531
          "011100100010100000110101" when "11000000", -- t[192] = 7481397
          "011100011111100100000011" when "11000001", -- t[193] = 7469315
          "011100011100101000000011" when "11000010", -- t[194] = 7457283
          "011100011001101100110110" when "11000011", -- t[195] = 7445302
          "011100010110110010011011" when "11000100", -- t[196] = 7433371
          "011100010011111000110010" when "11000101", -- t[197] = 7421490
          "011100010000111111111011" when "11000110", -- t[198] = 7409659
          "011100001110000111110101" when "11000111", -- t[199] = 7397877
          "011100001011010000011111" when "11001000", -- t[200] = 7386143
          "011100001000011001111011" when "11001001", -- t[201] = 7374459
          "011100000101100100000110" when "11001010", -- t[202] = 7362822
          "011100000010101111000001" when "11001011", -- t[203] = 7351233
          "011011111111111010101100" when "11001100", -- t[204] = 7339692
          "011011111101000111000110" when "11001101", -- t[205] = 7328198
          "011011111010010100001111" when "11001110", -- t[206] = 7316751
          "011011110111100010000110" when "11001111", -- t[207] = 7305350
          "011011110100110000101100" when "11010000", -- t[208] = 7293996
          "011011110010000000000000" when "11010001", -- t[209] = 7282688
          "011011101111010000000001" when "11010010", -- t[210] = 7271425
          "011011101100100000101111" when "11010011", -- t[211] = 7260207
          "011011101001110010001011" when "11010100", -- t[212] = 7249035
          "011011100111000100010011" when "11010101", -- t[213] = 7237907
          "011011100100010111001000" when "11010110", -- t[214] = 7226824
          "011011100001101010101001" when "11010111", -- t[215] = 7215785
          "011011011110111110110101" when "11011000", -- t[216] = 7204789
          "011011011100010011101101" when "11011001", -- t[217] = 7193837
          "011011011001101001010001" when "11011010", -- t[218] = 7182929
          "011011010110111111011111" when "11011011", -- t[219] = 7172063
          "011011010100010110011000" when "11011100", -- t[220] = 7161240
          "011011010001101101111100" when "11011101", -- t[221] = 7150460
          "011011001111000110001001" when "11011110", -- t[222] = 7139721
          "011011001100011111000000" when "11011111", -- t[223] = 7129024
          "011011001001111000100001" when "11100000", -- t[224] = 7118369
          "011011000111010010101100" when "11100001", -- t[225] = 7107756
          "011011000100101101011111" when "11100010", -- t[226] = 7097183
          "011011000010001000111011" when "11100011", -- t[227] = 7086651
          "011010111111100101000000" when "11100100", -- t[228] = 7076160
          "011010111101000001101100" when "11100101", -- t[229] = 7065708
          "011010111010011111000001" when "11100110", -- t[230] = 7055297
          "011010110111111100111110" when "11100111", -- t[231] = 7044926
          "011010110101011011100010" when "11101000", -- t[232] = 7034594
          "011010110010111010101101" when "11101001", -- t[233] = 7024301
          "011010110000011010011111" when "11101010", -- t[234] = 7014047
          "011010101101111010111000" when "11101011", -- t[235] = 7003832
          "011010101011011011111000" when "11101100", -- t[236] = 6993656
          "011010101000111101011110" when "11101101", -- t[237] = 6983518
          "011010100110011111101010" when "11101110", -- t[238] = 6973418
          "011010100100000010011011" when "11101111", -- t[239] = 6963355
          "011010100001100101110010" when "11110000", -- t[240] = 6953330
          "011010011111001001101111" when "11110001", -- t[241] = 6943343
          "011010011100101110010000" when "11110010", -- t[242] = 6933392
          "011010011010010011010111" when "11110011", -- t[243] = 6923479
          "011010010111111001000010" when "11110100", -- t[244] = 6913602
          "011010010101011111010001" when "11110101", -- t[245] = 6903761
          "011010010011000110000101" when "11110110", -- t[246] = 6893957
          "011010010000101101011100" when "11110111", -- t[247] = 6884188
          "011010001110010101011000" when "11111000", -- t[248] = 6874456
          "011010001011111101110110" when "11111001", -- t[249] = 6864758
          "011010001001100110111001" when "11111010", -- t[250] = 6855097
          "011010000111010000011110" when "11111011", -- t[251] = 6845470
          "011010000100111010100110" when "11111100", -- t[252] = 6835878
          "011010000010100101010001" when "11111101", -- t[253] = 6826321
          "011010000000010000011110" when "11111110", -- t[254] = 6816798
          "011001111101111100001101" when "11111111", -- t[255] = 6807309
          "------------------------" when others;

  r(23 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 12; mu_1 = 12; lambda_1 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20_t1_pow is
  port ( x : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_20_t1_pow is
  signal pp0 : std_logic_vector(10 downto 0);
  signal r0 : std_logic_vector(10 downto 0);
begin
  pp0(10) <= x(10);

  pp0(9) <= x(9);

  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(10 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 8; wO_1,1 = 16.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20_t1_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of fp_log_log_20_t1_t1 is
  signal x : std_logic_vector(7 downto 0);
begin
  x <= a;

  with x select
    r <= "1001110001010111" when "00000000", -- t[0] = 40023
         "1001101011010010" when "00000001", -- t[1] = 39634
         "1001100101010100" when "00000010", -- t[2] = 39252
         "1001011111011100" when "00000011", -- t[3] = 38876
         "1001011001101010" when "00000100", -- t[4] = 38506
         "1001010011111110" when "00000101", -- t[5] = 38142
         "1001001110011000" when "00000110", -- t[6] = 37784
         "1001001000111000" when "00000111", -- t[7] = 37432
         "1001000011011101" when "00001000", -- t[8] = 37085
         "1000111110001000" when "00001001", -- t[9] = 36744
         "1000111000111000" when "00001010", -- t[10] = 36408
         "1000110011101110" when "00001011", -- t[11] = 36078
         "1000101110101000" when "00001100", -- t[12] = 35752
         "1000101001101000" when "00001101", -- t[13] = 35432
         "1000100100101101" when "00001110", -- t[14] = 35117
         "1000011111110110" when "00001111", -- t[15] = 34806
         "1000011011000100" when "00010000", -- t[16] = 34500
         "1000010110010111" when "00010001", -- t[17] = 34199
         "1000010001101110" when "00010010", -- t[18] = 33902
         "1000001101001010" when "00010011", -- t[19] = 33610
         "1000001000101010" when "00010100", -- t[20] = 33322
         "1000000100001110" when "00010101", -- t[21] = 33038
         "0111111111110110" when "00010110", -- t[22] = 32758
         "0111111011100010" when "00010111", -- t[23] = 32482
         "0111110111010011" when "00011000", -- t[24] = 32211
         "0111110011000111" when "00011001", -- t[25] = 31943
         "0111101110111111" when "00011010", -- t[26] = 31679
         "0111101010111011" when "00011011", -- t[27] = 31419
         "0111100110111010" when "00011100", -- t[28] = 31162
         "0111100010111101" when "00011101", -- t[29] = 30909
         "0111011111000011" when "00011110", -- t[30] = 30659
         "0111011011001101" when "00011111", -- t[31] = 30413
         "0111010111011011" when "00100000", -- t[32] = 30171
         "0111010011101011" when "00100001", -- t[33] = 29931
         "0111001111111111" when "00100010", -- t[34] = 29695
         "0111001100010110" when "00100011", -- t[35] = 29462
         "0111001000110000" when "00100100", -- t[36] = 29232
         "0111000101001101" when "00100101", -- t[37] = 29005
         "0111000001101101" when "00100110", -- t[38] = 28781
         "0110111110010000" when "00100111", -- t[39] = 28560
         "0110111010110110" when "00101000", -- t[40] = 28342
         "0110110111011111" when "00101001", -- t[41] = 28127
         "0110110100001011" when "00101010", -- t[42] = 27915
         "0110110000111001" when "00101011", -- t[43] = 27705
         "0110101101101010" when "00101100", -- t[44] = 27498
         "0110101010011110" when "00101101", -- t[45] = 27294
         "0110100111010100" when "00101110", -- t[46] = 27092
         "0110100100001101" when "00101111", -- t[47] = 26893
         "0110100001001000" when "00110000", -- t[48] = 26696
         "0110011110000110" when "00110001", -- t[49] = 26502
         "0110011011000110" when "00110010", -- t[50] = 26310
         "0110011000001000" when "00110011", -- t[51] = 26120
         "0110010101001101" when "00110100", -- t[52] = 25933
         "0110010010010100" when "00110101", -- t[53] = 25748
         "0110001111011101" when "00110110", -- t[54] = 25565
         "0110001100101001" when "00110111", -- t[55] = 25385
         "0110001001110111" when "00111000", -- t[56] = 25207
         "0110000111000110" when "00111001", -- t[57] = 25030
         "0110000100011000" when "00111010", -- t[58] = 24856
         "0110000001101100" when "00111011", -- t[59] = 24684
         "0101111111000010" when "00111100", -- t[60] = 24514
         "0101111100011010" when "00111101", -- t[61] = 24346
         "0101111001110100" when "00111110", -- t[62] = 24180
         "0101110111010000" when "00111111", -- t[63] = 24016
         "0101110100101110" when "01000000", -- t[64] = 23854
         "0101110010001101" when "01000001", -- t[65] = 23693
         "0101101111101111" when "01000010", -- t[66] = 23535
         "0101101101010010" when "01000011", -- t[67] = 23378
         "0101101010110111" when "01000100", -- t[68] = 23223
         "0101101000011110" when "01000101", -- t[69] = 23070
         "0101100110000110" when "01000110", -- t[70] = 22918
         "0101100011110000" when "01000111", -- t[71] = 22768
         "0101100001011100" when "01001000", -- t[72] = 22620
         "0101011111001001" when "01001001", -- t[73] = 22473
         "0101011100111000" when "01001010", -- t[74] = 22328
         "0101011010101001" when "01001011", -- t[75] = 22185
         "0101011000011011" when "01001100", -- t[76] = 22043
         "0101010110001111" when "01001101", -- t[77] = 21903
         "0101010100000100" when "01001110", -- t[78] = 21764
         "0101010001111011" when "01001111", -- t[79] = 21627
         "0101001111110011" when "01010000", -- t[80] = 21491
         "0101001101101101" when "01010001", -- t[81] = 21357
         "0101001011101000" when "01010010", -- t[82] = 21224
         "0101001001100100" when "01010011", -- t[83] = 21092
         "0101000111100010" when "01010100", -- t[84] = 20962
         "0101000101100001" when "01010101", -- t[85] = 20833
         "0101000011100010" when "01010110", -- t[86] = 20706
         "0101000001100011" when "01010111", -- t[87] = 20579
         "0100111111100111" when "01011000", -- t[88] = 20455
         "0100111101101011" when "01011001", -- t[89] = 20331
         "0100111011110001" when "01011010", -- t[90] = 20209
         "0100111001111000" when "01011011", -- t[91] = 20088
         "0100111000000000" when "01011100", -- t[92] = 19968
         "0100110110001001" when "01011101", -- t[93] = 19849
         "0100110100010100" when "01011110", -- t[94] = 19732
         "0100110010011111" when "01011111", -- t[95] = 19615
         "0100110000101100" when "01100000", -- t[96] = 19500
         "0100101110111010" when "01100001", -- t[97] = 19386
         "0100101101001001" when "01100010", -- t[98] = 19273
         "0100101011011010" when "01100011", -- t[99] = 19162
         "0100101001101011" when "01100100", -- t[100] = 19051
         "0100100111111101" when "01100101", -- t[101] = 18941
         "0100100110010001" when "01100110", -- t[102] = 18833
         "0100100100100101" when "01100111", -- t[103] = 18725
         "0100100010111011" when "01101000", -- t[104] = 18619
         "0100100001010001" when "01101001", -- t[105] = 18513
         "0100011111101001" when "01101010", -- t[106] = 18409
         "0100011110000010" when "01101011", -- t[107] = 18306
         "0100011100011011" when "01101100", -- t[108] = 18203
         "0100011010110110" when "01101101", -- t[109] = 18102
         "0100011001010001" when "01101110", -- t[110] = 18001
         "0100010111101110" when "01101111", -- t[111] = 17902
         "0100010110001011" when "01110000", -- t[112] = 17803
         "0100010100101001" when "01110001", -- t[113] = 17705
         "0100010011001000" when "01110010", -- t[114] = 17608
         "0100010001101001" when "01110011", -- t[115] = 17513
         "0100010000001001" when "01110100", -- t[116] = 17417
         "0100001110101011" when "01110101", -- t[117] = 17323
         "0100001101001110" when "01110110", -- t[118] = 17230
         "0100001011110001" when "01110111", -- t[119] = 17137
         "0100001010010110" when "01111000", -- t[120] = 17046
         "0100001000111011" when "01111001", -- t[121] = 16955
         "0100000111100001" when "01111010", -- t[122] = 16865
         "0100000110001000" when "01111011", -- t[123] = 16776
         "0100000100101111" when "01111100", -- t[124] = 16687
         "0100000011011000" when "01111101", -- t[125] = 16600
         "0100000010000001" when "01111110", -- t[126] = 16513
         "0100000000101011" when "01111111", -- t[127] = 16427
         "0011111111010101" when "10000000", -- t[128] = 16341
         "0011111110000001" when "10000001", -- t[129] = 16257
         "0011111100101101" when "10000010", -- t[130] = 16173
         "0011111011011010" when "10000011", -- t[131] = 16090
         "0011111010000111" when "10000100", -- t[132] = 16007
         "0011111000110110" when "10000101", -- t[133] = 15926
         "0011110111100101" when "10000110", -- t[134] = 15845
         "0011110110010100" when "10000111", -- t[135] = 15764
         "0011110101000101" when "10001000", -- t[136] = 15685
         "0011110011110110" when "10001001", -- t[137] = 15606
         "0011110010101000" when "10001010", -- t[138] = 15528
         "0011110001011010" when "10001011", -- t[139] = 15450
         "0011110000001101" when "10001100", -- t[140] = 15373
         "0011101111000001" when "10001101", -- t[141] = 15297
         "0011101101110101" when "10001110", -- t[142] = 15221
         "0011101100101010" when "10001111", -- t[143] = 15146
         "0011101011100000" when "10010000", -- t[144] = 15072
         "0011101010010110" when "10010001", -- t[145] = 14998
         "0011101001001101" when "10010010", -- t[146] = 14925
         "0011101000000100" when "10010011", -- t[147] = 14852
         "0011100110111100" when "10010100", -- t[148] = 14780
         "0011100101110100" when "10010101", -- t[149] = 14708
         "0011100100101110" when "10010110", -- t[150] = 14638
         "0011100011100111" when "10010111", -- t[151] = 14567
         "0011100010100010" when "10011000", -- t[152] = 14498
         "0011100001011100" when "10011001", -- t[153] = 14428
         "0011100000011000" when "10011010", -- t[154] = 14360
         "0011011111010100" when "10011011", -- t[155] = 14292
         "0011011110010000" when "10011100", -- t[156] = 14224
         "0011011101001101" when "10011101", -- t[157] = 14157
         "0011011100001011" when "10011110", -- t[158] = 14091
         "0011011011001001" when "10011111", -- t[159] = 14025
         "0011011010000111" when "10100000", -- t[160] = 13959
         "0011011001000111" when "10100001", -- t[161] = 13895
         "0011011000000110" when "10100010", -- t[162] = 13830
         "0011010111000110" when "10100011", -- t[163] = 13766
         "0011010110000111" when "10100100", -- t[164] = 13703
         "0011010101001000" when "10100101", -- t[165] = 13640
         "0011010100001001" when "10100110", -- t[166] = 13577
         "0011010011001100" when "10100111", -- t[167] = 13516
         "0011010010001110" when "10101000", -- t[168] = 13454
         "0011010001010001" when "10101001", -- t[169] = 13393
         "0011010000010100" when "10101010", -- t[170] = 13332
         "0011001111011000" when "10101011", -- t[171] = 13272
         "0011001110011101" when "10101100", -- t[172] = 13213
         "0011001101100010" when "10101101", -- t[173] = 13154
         "0011001100100111" when "10101110", -- t[174] = 13095
         "0011001011101100" when "10101111", -- t[175] = 13036
         "0011001010110011" when "10110000", -- t[176] = 12979
         "0011001001111001" when "10110001", -- t[177] = 12921
         "0011001001000000" when "10110010", -- t[178] = 12864
         "0011001000001000" when "10110011", -- t[179] = 12808
         "0011000111001111" when "10110100", -- t[180] = 12751
         "0011000110011000" when "10110101", -- t[181] = 12696
         "0011000101100000" when "10110110", -- t[182] = 12640
         "0011000100101001" when "10110111", -- t[183] = 12585
         "0011000011110011" when "10111000", -- t[184] = 12531
         "0011000010111101" when "10111001", -- t[185] = 12477
         "0011000010000111" when "10111010", -- t[186] = 12423
         "0011000001010001" when "10111011", -- t[187] = 12369
         "0011000000011100" when "10111100", -- t[188] = 12316
         "0010111111101000" when "10111101", -- t[189] = 12264
         "0010111110110100" when "10111110", -- t[190] = 12212
         "0010111110000000" when "10111111", -- t[191] = 12160
         "0010111101001100" when "11000000", -- t[192] = 12108
         "0010111100011001" when "11000001", -- t[193] = 12057
         "0010111011100110" when "11000010", -- t[194] = 12006
         "0010111010110100" when "11000011", -- t[195] = 11956
         "0010111010000010" when "11000100", -- t[196] = 11906
         "0010111001010000" when "11000101", -- t[197] = 11856
         "0010111000011111" when "11000110", -- t[198] = 11807
         "0010110111101110" when "11000111", -- t[199] = 11758
         "0010110110111101" when "11001000", -- t[200] = 11709
         "0010110110001101" when "11001001", -- t[201] = 11661
         "0010110101011101" when "11001010", -- t[202] = 11613
         "0010110100101101" when "11001011", -- t[203] = 11565
         "0010110011111110" when "11001100", -- t[204] = 11518
         "0010110011001111" when "11001101", -- t[205] = 11471
         "0010110010100000" when "11001110", -- t[206] = 11424
         "0010110001110001" when "11001111", -- t[207] = 11377
         "0010110001000011" when "11010000", -- t[208] = 11331
         "0010110000010110" when "11010001", -- t[209] = 11286
         "0010101111101000" when "11010010", -- t[210] = 11240
         "0010101110111011" when "11010011", -- t[211] = 11195
         "0010101110001110" when "11010100", -- t[212] = 11150
         "0010101101100010" when "11010101", -- t[213] = 11106
         "0010101100110101" when "11010110", -- t[214] = 11061
         "0010101100001001" when "11010111", -- t[215] = 11017
         "0010101011011110" when "11011000", -- t[216] = 10974
         "0010101010110010" when "11011001", -- t[217] = 10930
         "0010101010000111" when "11011010", -- t[218] = 10887
         "0010101001011100" when "11011011", -- t[219] = 10844
         "0010101000110010" when "11011100", -- t[220] = 10802
         "0010101000000111" when "11011101", -- t[221] = 10759
         "0010100111011110" when "11011110", -- t[222] = 10718
         "0010100110110100" when "11011111", -- t[223] = 10676
         "0010100110001010" when "11100000", -- t[224] = 10634
         "0010100101100001" when "11100001", -- t[225] = 10593
         "0010100100111000" when "11100010", -- t[226] = 10552
         "0010100100010000" when "11100011", -- t[227] = 10512
         "0010100011100111" when "11100100", -- t[228] = 10471
         "0010100010111111" when "11100101", -- t[229] = 10431
         "0010100010010111" when "11100110", -- t[230] = 10391
         "0010100001110000" when "11100111", -- t[231] = 10352
         "0010100001001000" when "11101000", -- t[232] = 10312
         "0010100000100001" when "11101001", -- t[233] = 10273
         "0010011111111010" when "11101010", -- t[234] = 10234
         "0010011111010100" when "11101011", -- t[235] = 10196
         "0010011110101101" when "11101100", -- t[236] = 10157
         "0010011110000111" when "11101101", -- t[237] = 10119
         "0010011101100001" when "11101110", -- t[238] = 10081
         "0010011100111100" when "11101111", -- t[239] = 10044
         "0010011100010110" when "11110000", -- t[240] = 10006
         "0010011011110001" when "11110001", -- t[241] = 9969
         "0010011011001100" when "11110010", -- t[242] = 9932
         "0010011010100111" when "11110011", -- t[243] = 9895
         "0010011010000011" when "11110100", -- t[244] = 9859
         "0010011001011110" when "11110101", -- t[245] = 9822
         "0010011000111010" when "11110110", -- t[246] = 9786
         "0010011000010111" when "11110111", -- t[247] = 9751
         "0010010111110011" when "11111000", -- t[248] = 9715
         "0010010111001111" when "11111001", -- t[249] = 9679
         "0010010110101100" when "11111010", -- t[250] = 9644
         "0010010110001001" when "11111011", -- t[251] = 9609
         "0010010101100111" when "11111100", -- t[252] = 9575
         "0010010101000100" when "11111101", -- t[253] = 9540
         "0010010100100010" when "11111110", -- t[254] = 9506
         "0010010011111111" when "11111111", -- t[255] = 9471
         "----------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 8; beta_1 = 12; lambda_1 = 12;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 8; rho_1,1 = 0; sigma_1,1 = 12; wO_1,1 = 16.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         b : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(23 downto 0) );
end entity;

architecture arch of fp_log_log_20_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(10 downto 0);
  signal s      : std_logic_vector(11 downto 0);
  component fp_log_log_20_t1_pow is
    port ( x : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  signal a_1    : std_logic_vector(7 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(10 downto 0);
  signal k_1    : std_logic_vector(15 downto 0);
  signal r0_1   : std_logic_vector(28 downto 0);
  signal r_1    : std_logic_vector(23 downto 0);
  component fp_log_log_20_t1_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(15 downto 0) );
  end component;
begin
  sign <= not b(11);
  b0 <= b(10 downto 0) xor (10 downto 0 => sign);

  pow : fp_log_log_20_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(7 downto 0);
  sign_1 <= not s(11);
  s_1 <= s(10 downto 0) xor (10 downto 0 => sign_1);
  t_1 : fp_log_log_20_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(15 downto 0) <=
    r0_1(28 downto 13) xor (28 downto 13 => (not (sign xor sign_1)));
  r_1(23 downto 16) <= (23 downto 16 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 6; mu_2 = 12; lambda_2 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20_t2_pow is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_log_log_20_t2_pow is
  signal pp0 : std_logic_vector(10 downto 0);
  signal pp1 : std_logic_vector(10 downto 0);
  signal pp2 : std_logic_vector(10 downto 0);
  signal pp3 : std_logic_vector(10 downto 0);
  signal r0 : std_logic_vector(10 downto 0);
begin
  pp0(10) <= '0';
  pp1(10) <= '0';
  pp2(10) <= '0';
  pp3(10) <= '0';

  pp0(9) <= x(3) and x(4);
  pp1(9) <= x(4);
  pp2(9) <= '0';
  pp3(9) <= '0';

  pp0(8) <= x(2) and x(4);
  pp1(8) <= '0';
  pp2(8) <= '0';
  pp3(8) <= '0';

  pp0(7) <= x(1) and x(4);
  pp1(7) <= x(2) and x(3);
  pp2(7) <= x(3);
  pp3(7) <= '0';

  pp0(6) <= x(0) and x(4);
  pp1(6) <= x(1) and x(3);
  pp2(6) <= '0';
  pp3(6) <= '0';

  pp0(5) <= x(0) and x(3);
  pp1(5) <= x(1) and x(2);
  pp2(5) <= x(2);
  pp3(5) <= x(4);

  pp0(4) <= x(0) and x(2);
  pp1(4) <= x(3);
  pp2(4) <= '0';
  pp3(4) <= '0';

  pp0(3) <= x(0) and x(1);
  pp1(3) <= x(1);
  pp2(3) <= x(2);
  pp3(3) <= '0';

  pp0(2) <= x(0);
  pp1(2) <= x(1);
  pp2(2) <= '0';
  pp3(2) <= '0';

  pp0(1) <= '0';
  pp1(1) <= '0';
  pp2(1) <= '0';
  pp3(1) <= '0';

  pp0(0) <= '0';
  pp1(0) <= '0';
  pp2(0) <= '0';
  pp3(0) <= '0';

  r0 <= pp0 + pp1 + pp2 + pp3;
  r <= "1" & r0(10 downto 4);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 6; wO_2,1 = 7.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20_t2_t1 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of fp_log_log_20_t2_t1 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a;

  with x select
    r <= "1100000" when "000000", -- t[0] = 96
         "1011010" when "000001", -- t[1] = 90
         "1010100" when "000010", -- t[2] = 84
         "1001111" when "000011", -- t[3] = 79
         "1001010" when "000100", -- t[4] = 74
         "1000110" when "000101", -- t[5] = 70
         "1000010" when "000110", -- t[6] = 66
         "0111110" when "000111", -- t[7] = 62
         "0111011" when "001000", -- t[8] = 59
         "0111000" when "001001", -- t[9] = 56
         "0110101" when "001010", -- t[10] = 53
         "0110010" when "001011", -- t[11] = 50
         "0110000" when "001100", -- t[12] = 48
         "0101110" when "001101", -- t[13] = 46
         "0101100" when "001110", -- t[14] = 44
         "0101010" when "001111", -- t[15] = 42
         "0101000" when "010000", -- t[16] = 40
         "0100110" when "010001", -- t[17] = 38
         "0100100" when "010010", -- t[18] = 36
         "0100011" when "010011", -- t[19] = 35
         "0100001" when "010100", -- t[20] = 33
         "0100000" when "010101", -- t[21] = 32
         "0011111" when "010110", -- t[22] = 31
         "0011101" when "010111", -- t[23] = 29
         "0011100" when "011000", -- t[24] = 28
         "0011011" when "011001", -- t[25] = 27
         "0011010" when "011010", -- t[26] = 26
         "0011001" when "011011", -- t[27] = 25
         "0011000" when "011100", -- t[28] = 24
         "0010111" when "011101", -- t[29] = 23
         "0010111" when "011110", -- t[30] = 23
         "0010110" when "011111", -- t[31] = 22
         "0010101" when "100000", -- t[32] = 21
         "0010100" when "100001", -- t[33] = 20
         "0010100" when "100010", -- t[34] = 20
         "0010011" when "100011", -- t[35] = 19
         "0010010" when "100100", -- t[36] = 18
         "0010010" when "100101", -- t[37] = 18
         "0010001" when "100110", -- t[38] = 17
         "0010001" when "100111", -- t[39] = 17
         "0010000" when "101000", -- t[40] = 16
         "0010000" when "101001", -- t[41] = 16
         "0001111" when "101010", -- t[42] = 15
         "0001111" when "101011", -- t[43] = 15
         "0001110" when "101100", -- t[44] = 14
         "0001110" when "101101", -- t[45] = 14
         "0001101" when "101110", -- t[46] = 13
         "0001101" when "101111", -- t[47] = 13
         "0001101" when "110000", -- t[48] = 13
         "0001100" when "110001", -- t[49] = 12
         "0001100" when "110010", -- t[50] = 12
         "0001100" when "110011", -- t[51] = 12
         "0001011" when "110100", -- t[52] = 11
         "0001011" when "110101", -- t[53] = 11
         "0001011" when "110110", -- t[54] = 11
         "0001010" when "110111", -- t[55] = 10
         "0001010" when "111000", -- t[56] = 10
         "0001010" when "111001", -- t[57] = 10
         "0001010" when "111010", -- t[58] = 10
         "0001001" when "111011", -- t[59] = 9
         "0001001" when "111100", -- t[60] = 9
         "0001001" when "111101", -- t[61] = 9
         "0001001" when "111110", -- t[62] = 9
         "0001001" when "111111", -- t[63] = 9
         "-------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 6; beta_2 = 6; lambda_2 = 8;  m_2 = 1;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 6; rho_2,1 = 0; sigma_2,1 = 8; wO_2,1 = 7.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20_t2 is
  port ( a : in  std_logic_vector(5 downto 0);
         b : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(23 downto 0) );
end entity;

architecture arch of fp_log_log_20_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(4 downto 0);
  signal s      : std_logic_vector(7 downto 0);
  component fp_log_log_20_t2_pow is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  signal a_1    : std_logic_vector(5 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(6 downto 0);
  signal k_1    : std_logic_vector(6 downto 0);
  signal r0_1   : std_logic_vector(15 downto 0);
  signal r_1    : std_logic_vector(23 downto 0);
  component fp_log_log_20_t2_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;
begin
  sign <= not b(5);
  b0 <= b(4 downto 0) xor (4 downto 0 => sign);

  pow : fp_log_log_20_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(5 downto 0);
  sign_1 <= not s(7);
  s_1 <= s(6 downto 0) xor (6 downto 0 => sign_1);
  t_1 : fp_log_log_20_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(6 downto 0) <=
    r0_1(15 downto 9) xor (15 downto 9 => ((sign_1)));
  r_1(23 downto 7) <= (23 downto 7 => ((sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_20 is
  port ( x : in  std_logic_vector(19 downto 0);
         r : out std_logic_vector(23 downto 0) );
end entity;

architecture arch of fp_log_log_20 is
  signal a_0 : std_logic_vector(7 downto 0);
  signal r_0 : std_logic_vector(23 downto 0);
  component fp_log_log_20_t0 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(23 downto 0) );
  end component;

  signal a_1 : std_logic_vector(7 downto 0);
  signal b_1 : std_logic_vector(11 downto 0);
  signal r_1 : std_logic_vector(23 downto 0);
  component fp_log_log_20_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           b : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(23 downto 0) );
  end component;

  signal a_2 : std_logic_vector(5 downto 0);
  signal b_2 : std_logic_vector(5 downto 0);
  signal r_2 : std_logic_vector(23 downto 0);
  component fp_log_log_20_t2 is
    port ( a : in  std_logic_vector(5 downto 0);
           b : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(23 downto 0) );
  end component;

begin
  a_0 <= x(19 downto 12);
  t_0 : fp_log_log_20_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(19 downto 12);
  b_1 <= x(11 downto 0);
  t_1 : fp_log_log_20_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(19 downto 14);
  b_2 <= x(11 downto 6);
  t_2 : fp_log_log_20_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 21; wO = 21.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 8; beta = 13;
--   T_0 (ROM):     alpha_0 = 8; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 8; beta_1 = 13;
--   T_2 (PowMult): alpha_2 = 6; beta_2 = 8.
-- Guard bits: g = 3.
-- Command line: logfp 21 21 2   rom 8 0   pm 8 13  ah 13 13 13  1 0  8 13 0   pm 6 8  ah 8 16 12  1 1  6 8 0  3 4 8


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 8; beta_0 = 0; wO_0 = 25.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t0 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(24 downto 0) );
end entity;

architecture arch of fp_log_log_21_t0 is
  signal x0   : std_logic_vector(7 downto 0);
  signal r0   : std_logic_vector(24 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "1011000100100011101111111" when "00000000", -- t[0] = 23218047
          "1011000010001000001010110" when "00000001", -- t[1] = 23138390
          "1010111111101110000110000" when "00000010", -- t[2] = 23059504
          "1010111101010101100000001" when "00000011", -- t[3] = 22981377
          "1010111010111110011000001" when "00000100", -- t[4] = 22904001
          "1010111000101000101011010" when "00000101", -- t[5] = 22827354
          "1010110110010100011000100" when "00000110", -- t[6] = 22751428
          "1010110100000001011110101" when "00000111", -- t[7] = 22676213
          "1010110001101111111100101" when "00001000", -- t[8] = 22601701
          "1010101111011111110000000" when "00001001", -- t[9] = 22527872
          "1010101101010000111000000" when "00001010", -- t[10] = 22454720
          "1010101011000011010011011" when "00001011", -- t[11] = 22382235
          "1010101000110111000001000" when "00001100", -- t[12] = 22310408
          "1010100110101011111111000" when "00001101", -- t[13] = 22239224
          "1010100100100010001100100" when "00001110", -- t[14] = 22168676
          "1010100010011001101000001" when "00001111", -- t[15] = 22098753
          "1010100000010010010001010" when "00010000", -- t[16] = 22029450
          "1010011110001100000101111" when "00010001", -- t[17] = 21960751
          "1010011100000111000101010" when "00010010", -- t[18] = 21892650
          "1010011010000011001110011" when "00010011", -- t[19] = 21825139
          "1010011000000000100000010" when "00010100", -- t[20] = 21758210
          "1010010101111110111001011" when "00010101", -- t[21] = 21691851
          "1010010011111110011000111" when "00010110", -- t[22] = 21626055
          "1010010001111110111101111" when "00010111", -- t[23] = 21560815
          "1010010000000000100111101" when "00011000", -- t[24] = 21496125
          "1010001110000011010100011" when "00011001", -- t[25] = 21431971
          "1010001100000111000011101" when "00011010", -- t[26] = 21368349
          "1010001010001011110100100" when "00011011", -- t[27] = 21305252
          "1010001000010001100110010" when "00011100", -- t[28] = 21242674
          "1010000110011000010111100" when "00011101", -- t[29] = 21180604
          "1010000100100000000111011" when "00011110", -- t[30] = 21119035
          "1010000010101000110101011" when "00011111", -- t[31] = 21057963
          "1010000000110010100000110" when "00100000", -- t[32] = 20997382
          "1001111110111101001000000" when "00100001", -- t[33] = 20937280
          "1001111101001000101010110" when "00100010", -- t[34] = 20877654
          "1001111011010101001000010" when "00100011", -- t[35] = 20818498
          "1001111001100010011111110" when "00100100", -- t[36] = 20759806
          "1001110111110000110000010" when "00100101", -- t[37] = 20701570
          "1001110101111111111000111" when "00100110", -- t[38] = 20643783
          "1001110100001111111001010" when "00100111", -- t[39] = 20586442
          "1001110010100000110000110" when "00101000", -- t[40] = 20529542
          "1001110000110010011110001" when "00101001", -- t[41] = 20473073
          "1001101111000101000000111" when "00101010", -- t[42] = 20417031
          "1001101101011000011000011" when "00101011", -- t[43] = 20361411
          "1001101011101100100100010" when "00101100", -- t[44] = 20306210
          "1001101010000001100011011" when "00101101", -- t[45] = 20251419
          "1001101000010111010101001" when "00101110", -- t[46] = 20197033
          "1001100110101101111001001" when "00101111", -- t[47] = 20143049
          "1001100101000101001110110" when "00110000", -- t[48] = 20089462
          "1001100011011101010101001" when "00110001", -- t[49] = 20036265
          "1001100001110110001011101" when "00110010", -- t[50] = 19983453
          "1001100000001111110010000" when "00110011", -- t[51] = 19931024
          "1001011110101010000111100" when "00110100", -- t[52] = 19878972
          "1001011101000101001011011" when "00110101", -- t[53] = 19827291
          "1001011011100000111101010" when "00110110", -- t[54] = 19775978
          "1001011001111101011100100" when "00110111", -- t[55] = 19725028
          "1001011000011010101000110" when "00111000", -- t[56] = 19674438
          "1001010110111000100001010" when "00111001", -- t[57] = 19624202
          "1001010101010111000101011" when "00111010", -- t[58] = 19574315
          "1001010011110110010100111" when "00111011", -- t[59] = 19524775
          "1001010010010110001111010" when "00111100", -- t[60] = 19475578
          "1001010000110110110011110" when "00111101", -- t[61] = 19426718
          "1001001111011000000010000" when "00111110", -- t[62] = 19378192
          "1001001101111001111001100" when "00111111", -- t[63] = 19329996
          "1001001100011100011010000" when "01000000", -- t[64] = 19282128
          "1001001010111111100010101" when "01000001", -- t[65] = 19234581
          "1001001001100011010011010" when "01000010", -- t[66] = 19187354
          "1001001000000111101011010" when "01000011", -- t[67] = 19140442
          "1001000110101100101010010" when "01000100", -- t[68] = 19093842
          "1001000101010010001111110" when "01000101", -- t[69] = 19047550
          "1001000011111000011011011" when "01000110", -- t[70] = 19001563
          "1001000010011111001100101" when "01000111", -- t[71] = 18955877
          "1001000001000110100011010" when "01001000", -- t[72] = 18910490
          "1000111111101110011110101" when "01001001", -- t[73] = 18865397
          "1000111110010110111110100" when "01001010", -- t[74] = 18820596
          "1000111101000000000010010" when "01001011", -- t[75] = 18776082
          "1000111011101001101010000" when "01001100", -- t[76] = 18731856
          "1000111010010011110100110" when "01001101", -- t[77] = 18687910
          "1000111000111110100010011" when "01001110", -- t[78] = 18644243
          "1000110111101001110010100" when "01001111", -- t[79] = 18600852
          "1000110110010101100101000" when "01010000", -- t[80] = 18557736
          "1000110101000001111001000" when "01010001", -- t[81] = 18514888
          "1000110011101110101110100" when "01010010", -- t[82] = 18472308
          "1000110010011100000101001" when "01010011", -- t[83] = 18429993
          "1000110001001001111100100" when "01010100", -- t[84] = 18387940
          "1000101111111000010100001" when "01010101", -- t[85] = 18346145
          "1000101110100111001011111" when "01010110", -- t[86] = 18304607
          "1000101101010110100011010" when "01010111", -- t[87] = 18263322
          "1000101100000110011010001" when "01011000", -- t[88] = 18222289
          "1000101010110110110000000" when "01011001", -- t[89] = 18181504
          "1000101001100111100100100" when "01011010", -- t[90] = 18140964
          "1000101000011000110111100" when "01011011", -- t[91] = 18100668
          "1000100111001010101000110" when "01011100", -- t[92] = 18060614
          "1000100101111100110111101" when "01011101", -- t[93] = 18020797
          "1000100100101111100100001" when "01011110", -- t[94] = 17981217
          "1000100011100010101101110" when "01011111", -- t[95] = 17941870
          "1000100010010110010100100" when "01100000", -- t[96] = 17902756
          "1000100001001010010111101" when "01100001", -- t[97] = 17863869
          "1000011111111110110111010" when "01100010", -- t[98] = 17825210
          "1000011110110011110010111" when "01100011", -- t[99] = 17786775
          "1000011101101001001010100" when "01100100", -- t[100] = 17748564
          "1000011100011110111101011" when "01100101", -- t[101] = 17710571
          "1000011011010101001011101" when "01100110", -- t[102] = 17672797
          "1000011010001011110100111" when "01100111", -- t[103] = 17635239
          "1000011001000010111001000" when "01101000", -- t[104] = 17597896
          "1000010111111010010111100" when "01101001", -- t[105] = 17560764
          "1000010110110010010000001" when "01101010", -- t[106] = 17523841
          "1000010101101010100010110" when "01101011", -- t[107] = 17487126
          "1000010100100011001111010" when "01101100", -- t[108] = 17450618
          "1000010011011100010101001" when "01101101", -- t[109] = 17414313
          "1000010010010101110100010" when "01101110", -- t[110] = 17378210
          "1000010001001111101100100" when "01101111", -- t[111] = 17342308
          "1000010000001001111101100" when "01110000", -- t[112] = 17306604
          "1000001111000100100111000" when "01110001", -- t[113] = 17271096
          "1000001101111111101000110" when "01110010", -- t[114] = 17235782
          "1000001100111011000010101" when "01110011", -- t[115] = 17200661
          "1000001011110110110100100" when "01110100", -- t[116] = 17165732
          "1000001010110010111101111" when "01110101", -- t[117] = 17130991
          "1000001001101111011110110" when "01110110", -- t[118] = 17096438
          "1000001000101100010110110" when "01110111", -- t[119] = 17062070
          "1000000111101001100110000" when "01111000", -- t[120] = 17027888
          "1000000110100111001011111" when "01111001", -- t[121] = 16993887
          "1000000101100101001000011" when "01111010", -- t[122] = 16960067
          "1000000100100011011011010" when "01111011", -- t[123] = 16926426
          "1000000011100010000100100" when "01111100", -- t[124] = 16892964
          "1000000010100001000011101" when "01111101", -- t[125] = 16859677
          "1000000001100000011000100" when "01111110", -- t[126] = 16826564
          "1000000000100000000011001" when "01111111", -- t[127] = 16793625
          "0111111111100000000011001" when "10000000", -- t[128] = 16760857
          "0111111110100000011000011" when "10000001", -- t[129] = 16728259
          "0111111101100001000010101" when "10000010", -- t[130] = 16695829
          "0111111100100010000001110" when "10000011", -- t[131] = 16663566
          "0111111011100011010101101" when "10000100", -- t[132] = 16631469
          "0111111010100100111110000" when "10000101", -- t[133] = 16599536
          "0111111001100110111010101" when "10000110", -- t[134] = 16567765
          "0111111000101001001011100" when "10000111", -- t[135] = 16536156
          "0111110111101011110000011" when "10001000", -- t[136] = 16504707
          "0111110110101110101001001" when "10001001", -- t[137] = 16473417
          "0111110101110001110101011" when "10001010", -- t[138] = 16442283
          "0111110100110101010101001" when "10001011", -- t[139] = 16411305
          "0111110011111001001000011" when "10001100", -- t[140] = 16380483
          "0111110010111101001110101" when "10001101", -- t[141] = 16349813
          "0111110010000001100111111" when "10001110", -- t[142] = 16319295
          "0111110001000110010100000" when "10001111", -- t[143] = 16288928
          "0111110000001011010010111" when "10010000", -- t[144] = 16258711
          "0111101111010000100100010" when "10010001", -- t[145] = 16228642
          "0111101110010110001000000" when "10010010", -- t[146] = 16198720
          "0111101101011011111110000" when "10010011", -- t[147] = 16168944
          "0111101100100010000110000" when "10010100", -- t[148] = 16139312
          "0111101011101000100000000" when "10010101", -- t[149] = 16109824
          "0111101010101111001011110" when "10010110", -- t[150] = 16080478
          "0111101001110110001001001" when "10010111", -- t[151] = 16051273
          "0111101000111101011000001" when "10011000", -- t[152] = 16022209
          "0111101000000100111000011" when "10011001", -- t[153] = 15993283
          "0111100111001100101001111" when "10011010", -- t[154] = 15964495
          "0111100110010100101100011" when "10011011", -- t[155] = 15935843
          "0111100101011101000000000" when "10011100", -- t[156] = 15907328
          "0111100100100101100100010" when "10011101", -- t[157] = 15878946
          "0111100011101110011001010" when "10011110", -- t[158] = 15850698
          "0111100010110111011110111" when "10011111", -- t[159] = 15822583
          "0111100010000000110100111" when "10100000", -- t[160] = 15794599
          "0111100001001010011011001" when "10100001", -- t[161] = 15766745
          "0111100000010100010001101" when "10100010", -- t[162] = 15739021
          "0111011111011110011000000" when "10100011", -- t[163] = 15711424
          "0111011110101000101110100" when "10100100", -- t[164] = 15683956
          "0111011101110011010100101" when "10100101", -- t[165] = 15656613
          "0111011100111110001010100" when "10100110", -- t[166] = 15629396
          "0111011100001001001111111" when "10100111", -- t[167] = 15602303
          "0111011011010100100100110" when "10101000", -- t[168] = 15575334
          "0111011010100000001000111" when "10101001", -- t[169] = 15548487
          "0111011001101011111100001" when "10101010", -- t[170] = 15521761
          "0111011000110111111110100" when "10101011", -- t[171] = 15495156
          "0111011000000100010000000" when "10101100", -- t[172] = 15468672
          "0111010111010000110000001" when "10101101", -- t[173] = 15442305
          "0111010110011101011111001" when "10101110", -- t[174] = 15416057
          "0111010101101010011100110" when "10101111", -- t[175] = 15389926
          "0111010100110111101000111" when "10110000", -- t[176] = 15363911
          "0111010100000101000011011" when "10110001", -- t[177] = 15338011
          "0111010011010010101100010" when "10110010", -- t[178] = 15312226
          "0111010010100000100011010" when "10110011", -- t[179] = 15286554
          "0111010001101110101000011" when "10110100", -- t[180] = 15260995
          "0111010000111100111011100" when "10110101", -- t[181] = 15235548
          "0111010000001011011100101" when "10110110", -- t[182] = 15210213
          "0111001111011010001011011" when "10110111", -- t[183] = 15184987
          "0111001110101001000111111" when "10111000", -- t[184] = 15159871
          "0111001101111000010010000" when "10111001", -- t[185] = 15134864
          "0111001101000111101001101" when "10111010", -- t[186] = 15109965
          "0111001100010111001110100" when "10111011", -- t[187] = 15085172
          "0111001011100111000000111" when "10111100", -- t[188] = 15060487
          "0111001010110111000000011" when "10111101", -- t[189] = 15035907
          "0111001010000111001100111" when "10111110", -- t[190] = 15011431
          "0111001001010111100110100" when "10111111", -- t[191] = 14987060
          "0111001000101000001101000" when "11000000", -- t[192] = 14962792
          "0111000111111001000000011" when "11000001", -- t[193] = 14938627
          "0111000111001010000000100" when "11000010", -- t[194] = 14914564
          "0111000110011011001101010" when "11000011", -- t[195] = 14890602
          "0111000101101100100110100" when "11000100", -- t[196] = 14866740
          "0111000100111110001100010" when "11000101", -- t[197] = 14842978
          "0111000100001111111110100" when "11000110", -- t[198] = 14819316
          "0111000011100001111100111" when "11000111", -- t[199] = 14795751
          "0111000010110100000111101" when "11001000", -- t[200] = 14772285
          "0111000010000110011110011" when "11001001", -- t[201] = 14748915
          "0111000001011001000001010" when "11001010", -- t[202] = 14725642
          "0111000000101011110000001" when "11001011", -- t[203] = 14702465
          "0110111111111110101010110" when "11001100", -- t[204] = 14679382
          "0110111111010001110001010" when "11001101", -- t[205] = 14656394
          "0110111110100101000011100" when "11001110", -- t[206] = 14633500
          "0110111101111000100001011" when "11001111", -- t[207] = 14610699
          "0110111101001100001010110" when "11010000", -- t[208] = 14587990
          "0110111100011111111111110" when "11010001", -- t[209] = 14565374
          "0110111011110100000000000" when "11010010", -- t[210] = 14542848
          "0110111011001000001011101" when "11010011", -- t[211] = 14520413
          "0110111010011100100010100" when "11010100", -- t[212] = 14498068
          "0110111001110001000100101" when "11010101", -- t[213] = 14475813
          "0110111001000101110001110" when "11010110", -- t[214] = 14453646
          "0110111000011010101001111" when "11010111", -- t[215] = 14431567
          "0110110111101111101101001" when "11011000", -- t[216] = 14409577
          "0110110111000100111011001" when "11011001", -- t[217] = 14387673
          "0110110110011010010100000" when "11011010", -- t[218] = 14365856
          "0110110101101111110111100" when "11011011", -- t[219] = 14344124
          "0110110101000101100101110" when "11011100", -- t[220] = 14322478
          "0110110100011011011110101" when "11011101", -- t[221] = 14300917
          "0110110011110001100010000" when "11011110", -- t[222] = 14279440
          "0110110011000111101111111" when "11011111", -- t[223] = 14258047
          "0110110010011110001000001" when "11100000", -- t[224] = 14236737
          "0110110001110100101010101" when "11100001", -- t[225] = 14215509
          "0110110001001011010111100" when "11100010", -- t[226] = 14194364
          "0110110000100010001110100" when "11100011", -- t[227] = 14173300
          "0110101111111001001111101" when "11100100", -- t[228] = 14152317
          "0110101111010000011010111" when "11100101", -- t[229] = 14131415
          "0110101110100111110000001" when "11100110", -- t[230] = 14110593
          "0110101101111111001111010" when "11100111", -- t[231] = 14089850
          "0110101101010110111000010" when "11101000", -- t[232] = 14069186
          "0110101100101110101011000" when "11101001", -- t[233] = 14048600
          "0110101100000110100111101" when "11101010", -- t[234] = 14028093
          "0110101011011110101101111" when "11101011", -- t[235] = 14007663
          "0110101010110110111101110" when "11101100", -- t[236] = 13987310
          "0110101010001111010111010" when "11101101", -- t[237] = 13967034
          "0110101001100111111010001" when "11101110", -- t[238] = 13946833
          "0110101001000000100110101" when "11101111", -- t[239] = 13926709
          "0110101000011001011100011" when "11110000", -- t[240] = 13906659
          "0110100111110010011011100" when "11110001", -- t[241] = 13886684
          "0110100111001011100011111" when "11110010", -- t[242] = 13866783
          "0110100110100100110101100" when "11110011", -- t[243] = 13846956
          "0110100101111110010000010" when "11110100", -- t[244] = 13827202
          "0110100101010111110100001" when "11110101", -- t[245] = 13807521
          "0110100100110001100001000" when "11110110", -- t[246] = 13787912
          "0110100100001011010110111" when "11110111", -- t[247] = 13768375
          "0110100011100101010101110" when "11111000", -- t[248] = 13748910
          "0110100010111111011101011" when "11111001", -- t[249] = 13729515
          "0110100010011001101101111" when "11111010", -- t[250] = 13710191
          "0110100001110100000111010" when "11111011", -- t[251] = 13690938
          "0110100001001110101001010" when "11111100", -- t[252] = 13671754
          "0110100000101001010100000" when "11111101", -- t[253] = 13652640
          "0110100000000100000111010" when "11111110", -- t[254] = 13633594
          "0110011111011111000011001" when "11111111", -- t[255] = 13614617
          "-------------------------" when others;

  r(24 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 13; mu_1 = 13; lambda_1 = 13.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t1_pow is
  port ( x : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of fp_log_log_21_t1_pow is
  signal pp0 : std_logic_vector(11 downto 0);
  signal r0 : std_logic_vector(11 downto 0);
begin
  pp0(11) <= x(11);

  pp0(10) <= x(10);

  pp0(9) <= x(9);

  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(11 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 8; wO_1,1 = 17.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t1_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of fp_log_log_21_t1_t1 is
  signal x : std_logic_vector(7 downto 0);
begin
  x <= a;

  with x select
    r <= "10011100010101110" when "00000000", -- t[0] = 80046
         "10011010110100100" when "00000001", -- t[1] = 79268
         "10011001010100111" when "00000010", -- t[2] = 78503
         "10010111110110111" when "00000011", -- t[3] = 77751
         "10010110011010011" when "00000100", -- t[4] = 77011
         "10010100111111100" when "00000101", -- t[5] = 76284
         "10010011100110000" when "00000110", -- t[6] = 75568
         "10010010001101111" when "00000111", -- t[7] = 74863
         "10010000110111010" when "00001000", -- t[8] = 74170
         "10001111100010000" when "00001001", -- t[9] = 73488
         "10001110001110000" when "00001010", -- t[10] = 72816
         "10001100111011011" when "00001011", -- t[11] = 72155
         "10001011101010001" when "00001100", -- t[12] = 71505
         "10001010011010000" when "00001101", -- t[13] = 70864
         "10001001001011001" when "00001110", -- t[14] = 70233
         "10000111111101100" when "00001111", -- t[15] = 69612
         "10000110110001000" when "00010000", -- t[16] = 69000
         "10000101100101110" when "00010001", -- t[17] = 68398
         "10000100011011100" when "00010010", -- t[18] = 67804
         "10000011010010100" when "00010011", -- t[19] = 67220
         "10000010001010011" when "00010100", -- t[20] = 66643
         "10000001000011100" when "00010101", -- t[21] = 66076
         "01111111111101100" when "00010110", -- t[22] = 65516
         "01111110111000101" when "00010111", -- t[23] = 64965
         "01111101110100110" when "00011000", -- t[24] = 64422
         "01111100110001110" when "00011001", -- t[25] = 63886
         "01111011101111110" when "00011010", -- t[26] = 63358
         "01111010101110101" when "00011011", -- t[27] = 62837
         "01111001101110100" when "00011100", -- t[28] = 62324
         "01111000101111010" when "00011101", -- t[29] = 61818
         "01110111110000111" when "00011110", -- t[30] = 61319
         "01110110110011011" when "00011111", -- t[31] = 60827
         "01110101110110101" when "00100000", -- t[32] = 60341
         "01110100111010110" when "00100001", -- t[33] = 59862
         "01110011111111110" when "00100010", -- t[34] = 59390
         "01110011000101100" when "00100011", -- t[35] = 58924
         "01110010001100000" when "00100100", -- t[36] = 58464
         "01110001010011010" when "00100101", -- t[37] = 58010
         "01110000011011010" when "00100110", -- t[38] = 57562
         "01101111100100001" when "00100111", -- t[39] = 57121
         "01101110101101101" when "00101000", -- t[40] = 56685
         "01101101110111110" when "00101001", -- t[41] = 56254
         "01101101000010101" when "00101010", -- t[42] = 55829
         "01101100001110010" when "00101011", -- t[43] = 55410
         "01101011011010100" when "00101100", -- t[44] = 54996
         "01101010100111011" when "00101101", -- t[45] = 54587
         "01101001110101000" when "00101110", -- t[46] = 54184
         "01101001000011001" when "00101111", -- t[47] = 53785
         "01101000010010000" when "00110000", -- t[48] = 53392
         "01100111100001011" when "00110001", -- t[49] = 53003
         "01100110110001011" when "00110010", -- t[50] = 52619
         "01100110000010000" when "00110011", -- t[51] = 52240
         "01100101010011010" when "00110100", -- t[52] = 51866
         "01100100100101000" when "00110101", -- t[53] = 51496
         "01100011110111011" when "00110110", -- t[54] = 51131
         "01100011001010010" when "00110111", -- t[55] = 50770
         "01100010011101101" when "00111000", -- t[56] = 50413
         "01100001110001101" when "00111001", -- t[57] = 50061
         "01100001000110000" when "00111010", -- t[58] = 49712
         "01100000011011000" when "00111011", -- t[59] = 49368
         "01011111110000100" when "00111100", -- t[60] = 49028
         "01011111000110100" when "00111101", -- t[61] = 48692
         "01011110011101000" when "00111110", -- t[62] = 48360
         "01011101110100000" when "00111111", -- t[63] = 48032
         "01011101001011011" when "01000000", -- t[64] = 47707
         "01011100100011010" when "01000001", -- t[65] = 47386
         "01011011111011101" when "01000010", -- t[66] = 47069
         "01011011010100100" when "01000011", -- t[67] = 46756
         "01011010101101110" when "01000100", -- t[68] = 46446
         "01011010000111011" when "01000101", -- t[69] = 46139
         "01011001100001100" when "01000110", -- t[70] = 45836
         "01011000111100000" when "01000111", -- t[71] = 45536
         "01011000010111000" when "01001000", -- t[72] = 45240
         "01010111110010011" when "01001001", -- t[73] = 44947
         "01010111001110001" when "01001010", -- t[74] = 44657
         "01010110101010010" when "01001011", -- t[75] = 44370
         "01010110000110110" when "01001100", -- t[76] = 44086
         "01010101100011110" when "01001101", -- t[77] = 43806
         "01010101000001000" when "01001110", -- t[78] = 43528
         "01010100011110101" when "01001111", -- t[79] = 43253
         "01010011111100110" when "01010000", -- t[80] = 42982
         "01010011011011001" when "01010001", -- t[81] = 42713
         "01010010111001111" when "01010010", -- t[82] = 42447
         "01010010011001000" when "01010011", -- t[83] = 42184
         "01010001111000100" when "01010100", -- t[84] = 41924
         "01010001011000010" when "01010101", -- t[85] = 41666
         "01010000111000011" when "01010110", -- t[86] = 41411
         "01010000011000111" when "01010111", -- t[87] = 41159
         "01001111111001101" when "01011000", -- t[88] = 40909
         "01001111011010110" when "01011001", -- t[89] = 40662
         "01001110111100001" when "01011010", -- t[90] = 40417
         "01001110011101111" when "01011011", -- t[91] = 40175
         "01001101111111111" when "01011100", -- t[92] = 39935
         "01001101100010010" when "01011101", -- t[93] = 39698
         "01001101000100111" when "01011110", -- t[94] = 39463
         "01001100100111111" when "01011111", -- t[95] = 39231
         "01001100001011000" when "01100000", -- t[96] = 39000
         "01001011101110100" when "01100001", -- t[97] = 38772
         "01001011010010011" when "01100010", -- t[98] = 38547
         "01001010110110011" when "01100011", -- t[99] = 38323
         "01001010011010110" when "01100100", -- t[100] = 38102
         "01001001111111011" when "01100101", -- t[101] = 37883
         "01001001100100010" when "01100110", -- t[102] = 37666
         "01001001001001011" when "01100111", -- t[103] = 37451
         "01001000101110110" when "01101000", -- t[104] = 37238
         "01001000010100011" when "01101001", -- t[105] = 37027
         "01000111111010010" when "01101010", -- t[106] = 36818
         "01000111100000011" when "01101011", -- t[107] = 36611
         "01000111000110110" when "01101100", -- t[108] = 36406
         "01000110101101011" when "01101101", -- t[109] = 36203
         "01000110010100010" when "01101110", -- t[110] = 36002
         "01000101111011011" when "01101111", -- t[111] = 35803
         "01000101100010110" when "01110000", -- t[112] = 35606
         "01000101001010011" when "01110001", -- t[113] = 35411
         "01000100110010001" when "01110010", -- t[114] = 35217
         "01000100011010001" when "01110011", -- t[115] = 35025
         "01000100000010011" when "01110100", -- t[116] = 34835
         "01000011101010111" when "01110101", -- t[117] = 34647
         "01000011010011100" when "01110110", -- t[118] = 34460
         "01000010111100011" when "01110111", -- t[119] = 34275
         "01000010100101100" when "01111000", -- t[120] = 34092
         "01000010001110110" when "01111001", -- t[121] = 33910
         "01000001111000010" when "01111010", -- t[122] = 33730
         "01000001100010000" when "01111011", -- t[123] = 33552
         "01000001001011111" when "01111100", -- t[124] = 33375
         "01000000110101111" when "01111101", -- t[125] = 33199
         "01000000100000010" when "01111110", -- t[126] = 33026
         "01000000001010110" when "01111111", -- t[127] = 32854
         "00111111110101011" when "10000000", -- t[128] = 32683
         "00111111100000010" when "10000001", -- t[129] = 32514
         "00111111001011010" when "10000010", -- t[130] = 32346
         "00111110110110100" when "10000011", -- t[131] = 32180
         "00111110100001111" when "10000100", -- t[132] = 32015
         "00111110001101100" when "10000101", -- t[133] = 31852
         "00111101111001010" when "10000110", -- t[134] = 31690
         "00111101100101001" when "10000111", -- t[135] = 31529
         "00111101010001010" when "10001000", -- t[136] = 31370
         "00111100111101100" when "10001001", -- t[137] = 31212
         "00111100101001111" when "10001010", -- t[138] = 31055
         "00111100010110100" when "10001011", -- t[139] = 30900
         "00111100000011010" when "10001100", -- t[140] = 30746
         "00111011110000001" when "10001101", -- t[141] = 30593
         "00111011011101010" when "10001110", -- t[142] = 30442
         "00111011001010100" when "10001111", -- t[143] = 30292
         "00111010110111111" when "10010000", -- t[144] = 30143
         "00111010100101011" when "10010001", -- t[145] = 29995
         "00111010010011001" when "10010010", -- t[146] = 29849
         "00111010000001000" when "10010011", -- t[147] = 29704
         "00111001101111000" when "10010100", -- t[148] = 29560
         "00111001011101001" when "10010101", -- t[149] = 29417
         "00111001001011011" when "10010110", -- t[150] = 29275
         "00111000111001111" when "10010111", -- t[151] = 29135
         "00111000101000011" when "10011000", -- t[152] = 28995
         "00111000010111001" when "10011001", -- t[153] = 28857
         "00111000000110000" when "10011010", -- t[154] = 28720
         "00110111110100111" when "10011011", -- t[155] = 28583
         "00110111100100000" when "10011100", -- t[156] = 28448
         "00110111010011010" when "10011101", -- t[157] = 28314
         "00110111000010110" when "10011110", -- t[158] = 28182
         "00110110110010010" when "10011111", -- t[159] = 28050
         "00110110100001111" when "10100000", -- t[160] = 27919
         "00110110010001101" when "10100001", -- t[161] = 27789
         "00110110000001100" when "10100010", -- t[162] = 27660
         "00110101110001100" when "10100011", -- t[163] = 27532
         "00110101100001110" when "10100100", -- t[164] = 27406
         "00110101010010000" when "10100101", -- t[165] = 27280
         "00110101000010011" when "10100110", -- t[166] = 27155
         "00110100110010111" when "10100111", -- t[167] = 27031
         "00110100100011100" when "10101000", -- t[168] = 26908
         "00110100010100010" when "10101001", -- t[169] = 26786
         "00110100000101001" when "10101010", -- t[170] = 26665
         "00110011110110001" when "10101011", -- t[171] = 26545
         "00110011100111001" when "10101100", -- t[172] = 26425
         "00110011011000011" when "10101101", -- t[173] = 26307
         "00110011001001110" when "10101110", -- t[174] = 26190
         "00110010111011001" when "10101111", -- t[175] = 26073
         "00110010101100101" when "10110000", -- t[176] = 25957
         "00110010011110010" when "10110001", -- t[177] = 25842
         "00110010010000000" when "10110010", -- t[178] = 25728
         "00110010000001111" when "10110011", -- t[179] = 25615
         "00110001110011111" when "10110100", -- t[180] = 25503
         "00110001100101111" when "10110101", -- t[181] = 25391
         "00110001011000001" when "10110110", -- t[182] = 25281
         "00110001001010011" when "10110111", -- t[183] = 25171
         "00110000111100101" when "10111000", -- t[184] = 25061
         "00110000101111001" when "10111001", -- t[185] = 24953
         "00110000100001110" when "10111010", -- t[186] = 24846
         "00110000010100011" when "10111011", -- t[187] = 24739
         "00110000000111001" when "10111100", -- t[188] = 24633
         "00101111111010000" when "10111101", -- t[189] = 24528
         "00101111101100111" when "10111110", -- t[190] = 24423
         "00101111011111111" when "10111111", -- t[191] = 24319
         "00101111010011000" when "11000000", -- t[192] = 24216
         "00101111000110010" when "11000001", -- t[193] = 24114
         "00101110111001101" when "11000010", -- t[194] = 24013
         "00101110101101000" when "11000011", -- t[195] = 23912
         "00101110100000100" when "11000100", -- t[196] = 23812
         "00101110010100000" when "11000101", -- t[197] = 23712
         "00101110000111101" when "11000110", -- t[198] = 23613
         "00101101111011011" when "11000111", -- t[199] = 23515
         "00101101101111010" when "11001000", -- t[200] = 23418
         "00101101100011001" when "11001001", -- t[201] = 23321
         "00101101010111001" when "11001010", -- t[202] = 23225
         "00101101001011010" when "11001011", -- t[203] = 23130
         "00101100111111011" when "11001100", -- t[204] = 23035
         "00101100110011101" when "11001101", -- t[205] = 22941
         "00101100101000000" when "11001110", -- t[206] = 22848
         "00101100011100011" when "11001111", -- t[207] = 22755
         "00101100010000111" when "11010000", -- t[208] = 22663
         "00101100000101011" when "11010001", -- t[209] = 22571
         "00101011111010000" when "11010010", -- t[210] = 22480
         "00101011101110110" when "11010011", -- t[211] = 22390
         "00101011100011100" when "11010100", -- t[212] = 22300
         "00101011011000011" when "11010101", -- t[213] = 22211
         "00101011001101010" when "11010110", -- t[214] = 22122
         "00101011000010011" when "11010111", -- t[215] = 22035
         "00101010110111011" when "11011000", -- t[216] = 21947
         "00101010101100100" when "11011001", -- t[217] = 21860
         "00101010100001110" when "11011010", -- t[218] = 21774
         "00101010010111001" when "11011011", -- t[219] = 21689
         "00101010001100100" when "11011100", -- t[220] = 21604
         "00101010000001111" when "11011101", -- t[221] = 21519
         "00101001110111011" when "11011110", -- t[222] = 21435
         "00101001101101000" when "11011111", -- t[223] = 21352
         "00101001100010101" when "11100000", -- t[224] = 21269
         "00101001011000010" when "11100001", -- t[225] = 21186
         "00101001001110001" when "11100010", -- t[226] = 21105
         "00101001000011111" when "11100011", -- t[227] = 21023
         "00101000111001111" when "11100100", -- t[228] = 20943
         "00101000101111110" when "11100101", -- t[229] = 20862
         "00101000100101111" when "11100110", -- t[230] = 20783
         "00101000011011111" when "11100111", -- t[231] = 20703
         "00101000010010001" when "11101000", -- t[232] = 20625
         "00101000001000010" when "11101001", -- t[233] = 20546
         "00100111111110101" when "11101010", -- t[234] = 20469
         "00100111110100111" when "11101011", -- t[235] = 20391
         "00100111101011011" when "11101100", -- t[236] = 20315
         "00100111100001110" when "11101101", -- t[237] = 20238
         "00100111011000011" when "11101110", -- t[238] = 20163
         "00100111001110111" when "11101111", -- t[239] = 20087
         "00100111000101100" when "11110000", -- t[240] = 20012
         "00100110111100010" when "11110001", -- t[241] = 19938
         "00100110110011000" when "11110010", -- t[242] = 19864
         "00100110101001111" when "11110011", -- t[243] = 19791
         "00100110100000101" when "11110100", -- t[244] = 19717
         "00100110010111101" when "11110101", -- t[245] = 19645
         "00100110001110101" when "11110110", -- t[246] = 19573
         "00100110000101101" when "11110111", -- t[247] = 19501
         "00100101111100110" when "11111000", -- t[248] = 19430
         "00100101110011111" when "11111001", -- t[249] = 19359
         "00100101101011001" when "11111010", -- t[250] = 19289
         "00100101100010011" when "11111011", -- t[251] = 19219
         "00100101011001101" when "11111100", -- t[252] = 19149
         "00100101010001000" when "11111101", -- t[253] = 19080
         "00100101001000011" when "11111110", -- t[254] = 19011
         "00100100111111111" when "11111111", -- t[255] = 18943
         "-----------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 8; beta_1 = 13; lambda_1 = 13;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 8; rho_1,1 = 0; sigma_1,1 = 13; wO_1,1 = 17.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         b : in  std_logic_vector(12 downto 0);
         r : out std_logic_vector(24 downto 0) );
end entity;

architecture arch of fp_log_log_21_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(11 downto 0);
  signal s      : std_logic_vector(12 downto 0);
  component fp_log_log_21_t1_pow is
    port ( x : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  signal a_1    : std_logic_vector(7 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(11 downto 0);
  signal k_1    : std_logic_vector(16 downto 0);
  signal r0_1   : std_logic_vector(30 downto 0);
  signal r_1    : std_logic_vector(24 downto 0);
  component fp_log_log_21_t1_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(16 downto 0) );
  end component;
begin
  sign <= not b(12);
  b0 <= b(11 downto 0) xor (11 downto 0 => sign);

  pow : fp_log_log_21_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(7 downto 0);
  sign_1 <= not s(12);
  s_1 <= s(11 downto 0) xor (11 downto 0 => sign_1);
  t_1 : fp_log_log_21_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(16 downto 0) <=
    r0_1(30 downto 14) xor (30 downto 14 => (not (sign xor sign_1)));
  r_1(24 downto 17) <= (24 downto 17 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 8; mu_2 = 16; lambda_2 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t2_pow is
  port ( x : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_21_t2_pow is
  signal pp0 : std_logic_vector(14 downto 0);
  signal pp1 : std_logic_vector(14 downto 0);
  signal pp2 : std_logic_vector(14 downto 0);
  signal pp3 : std_logic_vector(14 downto 0);
  signal pp4 : std_logic_vector(14 downto 0);
  signal r0 : std_logic_vector(14 downto 0);
begin
  pp0(14) <= '0';
  pp1(14) <= '0';
  pp2(14) <= '0';
  pp3(14) <= '0';
  pp4(14) <= '0';

  pp0(13) <= x(5) and x(6);
  pp1(13) <= x(6);
  pp2(13) <= '0';
  pp3(13) <= '0';
  pp4(13) <= '0';

  pp0(12) <= x(4) and x(6);
  pp1(12) <= '0';
  pp2(12) <= '0';
  pp3(12) <= '0';
  pp4(12) <= '0';

  pp0(11) <= x(3) and x(6);
  pp1(11) <= x(4) and x(5);
  pp2(11) <= x(5);
  pp3(11) <= '0';
  pp4(11) <= '0';

  pp0(10) <= x(2) and x(6);
  pp1(10) <= x(3) and x(5);
  pp2(10) <= '0';
  pp3(10) <= '0';
  pp4(10) <= '0';

  pp0(9) <= x(1) and x(6);
  pp1(9) <= x(2) and x(5);
  pp2(9) <= x(3) and x(4);
  pp3(9) <= x(4);
  pp4(9) <= '0';

  pp0(8) <= x(0) and x(6);
  pp1(8) <= x(1) and x(5);
  pp2(8) <= x(2) and x(4);
  pp3(8) <= '0';
  pp4(8) <= '0';

  pp0(7) <= x(0) and x(5);
  pp1(7) <= x(1) and x(4);
  pp2(7) <= x(2) and x(3);
  pp3(7) <= x(3);
  pp4(7) <= x(6);

  pp0(6) <= x(0) and x(4);
  pp1(6) <= x(1) and x(3);
  pp2(6) <= x(5);
  pp3(6) <= '0';
  pp4(6) <= '0';

  pp0(5) <= x(0) and x(3);
  pp1(5) <= x(1) and x(2);
  pp2(5) <= x(2);
  pp3(5) <= x(4);
  pp4(5) <= '0';

  pp0(4) <= x(0) and x(2);
  pp1(4) <= x(3);
  pp2(4) <= '0';
  pp3(4) <= '0';
  pp4(4) <= '0';

  pp0(3) <= x(0) and x(1);
  pp1(3) <= x(1);
  pp2(3) <= x(2);
  pp3(3) <= '0';
  pp4(3) <= '0';

  pp0(2) <= x(0);
  pp1(2) <= x(1);
  pp2(2) <= '0';
  pp3(2) <= '0';
  pp4(2) <= '0';

  pp0(1) <= '0';
  pp1(1) <= '0';
  pp2(1) <= '0';
  pp3(1) <= '0';
  pp4(1) <= '0';

  pp0(0) <= '0';
  pp1(0) <= '0';
  pp2(0) <= '0';
  pp3(0) <= '0';
  pp4(0) <= '0';

  r0 <= pp0 + pp1 + pp2 + pp3 + pp4;
  r <= "1" & r0(14 downto 4);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 6; wO_2,1 = 8.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t2_t1 is
  port ( a : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of fp_log_log_21_t2_t1 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a;

  with x select
    r <= "10111111" when "000000", -- t[0] = 191
         "10110011" when "000001", -- t[1] = 179
         "10101000" when "000010", -- t[2] = 168
         "10011110" when "000011", -- t[3] = 158
         "10010100" when "000100", -- t[4] = 148
         "10001100" when "000101", -- t[5] = 140
         "10000100" when "000110", -- t[6] = 132
         "01111101" when "000111", -- t[7] = 125
         "01110110" when "001000", -- t[8] = 118
         "01110000" when "001001", -- t[9] = 112
         "01101010" when "001010", -- t[10] = 106
         "01100101" when "001011", -- t[11] = 101
         "01100000" when "001100", -- t[12] = 96
         "01011011" when "001101", -- t[13] = 91
         "01010111" when "001110", -- t[14] = 87
         "01010011" when "001111", -- t[15] = 83
         "01001111" when "010000", -- t[16] = 79
         "01001100" when "010001", -- t[17] = 76
         "01001000" when "010010", -- t[18] = 72
         "01000101" when "010011", -- t[19] = 69
         "01000010" when "010100", -- t[20] = 66
         "01000000" when "010101", -- t[21] = 64
         "00111101" when "010110", -- t[22] = 61
         "00111011" when "010111", -- t[23] = 59
         "00111000" when "011000", -- t[24] = 56
         "00110110" when "011001", -- t[25] = 54
         "00110100" when "011010", -- t[26] = 52
         "00110010" when "011011", -- t[27] = 50
         "00110000" when "011100", -- t[28] = 48
         "00101111" when "011101", -- t[29] = 47
         "00101101" when "011110", -- t[30] = 45
         "00101011" when "011111", -- t[31] = 43
         "00101010" when "100000", -- t[32] = 42
         "00101001" when "100001", -- t[33] = 41
         "00100111" when "100010", -- t[34] = 39
         "00100110" when "100011", -- t[35] = 38
         "00100101" when "100100", -- t[36] = 37
         "00100011" when "100101", -- t[37] = 35
         "00100010" when "100110", -- t[38] = 34
         "00100001" when "100111", -- t[39] = 33
         "00100000" when "101000", -- t[40] = 32
         "00011111" when "101001", -- t[41] = 31
         "00011110" when "101010", -- t[42] = 30
         "00011101" when "101011", -- t[43] = 29
         "00011101" when "101100", -- t[44] = 29
         "00011100" when "101101", -- t[45] = 28
         "00011011" when "101110", -- t[46] = 27
         "00011010" when "101111", -- t[47] = 26
         "00011001" when "110000", -- t[48] = 25
         "00011001" when "110001", -- t[49] = 25
         "00011000" when "110010", -- t[50] = 24
         "00010111" when "110011", -- t[51] = 23
         "00010111" when "110100", -- t[52] = 23
         "00010110" when "110101", -- t[53] = 22
         "00010110" when "110110", -- t[54] = 22
         "00010101" when "110111", -- t[55] = 21
         "00010100" when "111000", -- t[56] = 20
         "00010100" when "111001", -- t[57] = 20
         "00010011" when "111010", -- t[58] = 19
         "00010011" when "111011", -- t[59] = 19
         "00010010" when "111100", -- t[60] = 18
         "00010010" when "111101", -- t[61] = 18
         "00010010" when "111110", -- t[62] = 18
         "00010001" when "111111", -- t[63] = 17
         "--------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_2.
-- Decomposition:
--   alpha_2,2 = 3; sigma'_2,2 = 3; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t2_t2 is
  port ( a : in  std_logic_vector(2 downto 0);
         s : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of fp_log_log_21_t2_t2 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0" when "000000", -- t[0] = 0
         "0" when "000001", -- t[1] = 0
         "0" when "000010", -- t[2] = 0
         "0" when "000011", -- t[3] = 0
         "0" when "000100", -- t[4] = 0
         "0" when "000101", -- t[5] = 0
         "0" when "000110", -- t[6] = 0
         "0" when "000111", -- t[7] = 0
         "0" when "001000", -- t[8] = 0
         "0" when "001001", -- t[9] = 0
         "0" when "001010", -- t[10] = 0
         "0" when "001011", -- t[11] = 0
         "0" when "001100", -- t[12] = 0
         "0" when "001101", -- t[13] = 0
         "0" when "001110", -- t[14] = 0
         "0" when "001111", -- t[15] = 0
         "0" when "010000", -- t[16] = 0
         "0" when "010001", -- t[17] = 0
         "0" when "010010", -- t[18] = 0
         "0" when "010011", -- t[19] = 0
         "0" when "010100", -- t[20] = 0
         "0" when "010101", -- t[21] = 0
         "0" when "010110", -- t[22] = 0
         "0" when "010111", -- t[23] = 0
         "0" when "011000", -- t[24] = 0
         "0" when "011001", -- t[25] = 0
         "0" when "011010", -- t[26] = 0
         "0" when "011011", -- t[27] = 0
         "0" when "011100", -- t[28] = 0
         "0" when "011101", -- t[29] = 0
         "0" when "011110", -- t[30] = 0
         "0" when "011111", -- t[31] = 0
         "0" when "100000", -- t[32] = 0
         "0" when "100001", -- t[33] = 0
         "0" when "100010", -- t[34] = 0
         "0" when "100011", -- t[35] = 0
         "0" when "100100", -- t[36] = 0
         "0" when "100101", -- t[37] = 0
         "0" when "100110", -- t[38] = 0
         "0" when "100111", -- t[39] = 0
         "0" when "101000", -- t[40] = 0
         "0" when "101001", -- t[41] = 0
         "0" when "101010", -- t[42] = 0
         "0" when "101011", -- t[43] = 0
         "0" when "101100", -- t[44] = 0
         "0" when "101101", -- t[45] = 0
         "0" when "101110", -- t[46] = 0
         "0" when "101111", -- t[47] = 0
         "0" when "110000", -- t[48] = 0
         "0" when "110001", -- t[49] = 0
         "0" when "110010", -- t[50] = 0
         "0" when "110011", -- t[51] = 0
         "0" when "110100", -- t[52] = 0
         "0" when "110101", -- t[53] = 0
         "0" when "110110", -- t[54] = 0
         "0" when "110111", -- t[55] = 0
         "0" when "111000", -- t[56] = 0
         "0" when "111001", -- t[57] = 0
         "0" when "111010", -- t[58] = 0
         "0" when "111011", -- t[59] = 0
         "0" when "111100", -- t[60] = 0
         "0" when "111101", -- t[61] = 0
         "0" when "111110", -- t[62] = 0
         "0" when "111111", -- t[63] = 0
         "-" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 6; beta_2 = 8; lambda_2 = 12;  m_2 = 2;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 6; rho_2,1 = 0; sigma_2,1 = 8; wO_2,1 = 8;
--   Q_2,2 (ROM):  alpha_2,2 = 3; rho_2,2 = 8; sigma_2,2 = 4; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21_t2 is
  port ( a : in  std_logic_vector(5 downto 0);
         b : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(24 downto 0) );
end entity;

architecture arch of fp_log_log_21_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(6 downto 0);
  signal s      : std_logic_vector(11 downto 0);
  component fp_log_log_21_t2_pow is
    port ( x : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  signal a_1    : std_logic_vector(5 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(6 downto 0);
  signal k_1    : std_logic_vector(7 downto 0);
  signal r0_1   : std_logic_vector(16 downto 0);
  signal r_1    : std_logic_vector(24 downto 0);
  component fp_log_log_21_t2_t1 is
    port ( a : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  signal a_2    : std_logic_vector(2 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(2 downto 0);
  signal r0_2   : std_logic_vector(0 downto 0);
  signal r_2    : std_logic_vector(24 downto 0);
  component fp_log_log_21_t2_t2 is
    port ( a : in  std_logic_vector(2 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;
begin
  sign <= not b(7);
  b0 <= b(6 downto 0) xor (6 downto 0 => sign);

  pow : fp_log_log_21_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(5 downto 0);
  sign_1 <= not s(11);
  s_1 <= s(10 downto 4) xor (10 downto 4 => sign_1);
  t_1 : fp_log_log_21_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(7 downto 0) <=
    r0_1(16 downto 9) xor (16 downto 9 => ((sign_1)));
  r_1(24 downto 8) <= (24 downto 8 => ((sign_1)));

  a_2 <= a(5 downto 3);
  sign_2 <= not s(3);
  s_2 <= s(2 downto 0) xor (2 downto 0 => sign_2);
  t_2 : fp_log_log_21_t2_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(0 downto 0) <=
    r0_2 xor (0 downto 0 => ((sign_2)));
  r_2(24 downto 1) <= (24 downto 1 => ((sign_2)));

  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_21 is
  port ( x : in  std_logic_vector(20 downto 0);
         r : out std_logic_vector(24 downto 0) );
end entity;

architecture arch of fp_log_log_21 is
  signal a_0 : std_logic_vector(7 downto 0);
  signal r_0 : std_logic_vector(24 downto 0);
  component fp_log_log_21_t0 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(24 downto 0) );
  end component;

  signal a_1 : std_logic_vector(7 downto 0);
  signal b_1 : std_logic_vector(12 downto 0);
  signal r_1 : std_logic_vector(24 downto 0);
  component fp_log_log_21_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           b : in  std_logic_vector(12 downto 0);
           r : out std_logic_vector(24 downto 0) );
  end component;

  signal a_2 : std_logic_vector(5 downto 0);
  signal b_2 : std_logic_vector(7 downto 0);
  signal r_2 : std_logic_vector(24 downto 0);
  component fp_log_log_21_t2 is
    port ( a : in  std_logic_vector(5 downto 0);
           b : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(24 downto 0) );
  end component;

begin
  a_0 <= x(20 downto 13);
  t_0 : fp_log_log_21_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(20 downto 13);
  b_1 <= x(12 downto 0);
  t_1 : fp_log_log_21_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(20 downto 15);
  b_2 <= x(12 downto 5);
  t_2 : fp_log_log_21_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 22; wO = 22.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 8; beta = 14;
--   T_0 (ROM):     alpha_0 = 8; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 8; beta_1 = 14;
--   T_2 (PowMult): alpha_2 = 7; beta_2 = 8.
-- Guard bits: g = 3.
-- Command line: logfp 22 22 2   rom 8 0   pm 8 14  ah 14 14 14  1 0  8 14 0   pm 7 8  ah 8 16 12  1 1  7 8 0  3 4 8


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 8; beta_0 = 0; wO_0 = 26.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t0 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(25 downto 0) );
end entity;

architecture arch of fp_log_log_22_t0 is
  signal x0   : std_logic_vector(7 downto 0);
  signal r0   : std_logic_vector(25 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110001001000111011110101" when "00000000", -- t[0] = 46436085
          "10110000100010000010100011" when "00000001", -- t[1] = 46276771
          "10101111111011100001011101" when "00000010", -- t[2] = 46119005
          "10101111010101010111111110" when "00000011", -- t[3] = 45962750
          "10101110101111100101111001" when "00000100", -- t[4] = 45807993
          "10101110001010001010101010" when "00000101", -- t[5] = 45654698
          "10101101100101000110000100" when "00000110", -- t[6] = 45502852
          "10101101000000010111100110" when "00000111", -- t[7] = 45352422
          "10101100011011111111000010" when "00001000", -- t[8] = 45203394
          "10101011110111111011111000" when "00001001", -- t[9] = 45055736
          "10101011010100001101111101" when "00001010", -- t[10] = 44909437
          "10101010110000110100110001" when "00001011", -- t[11] = 44764465
          "10101010001101110000001001" when "00001100", -- t[12] = 44620809
          "10101001101010111111101001" when "00001101", -- t[13] = 44478441
          "10101001001000100011000011" when "00001110", -- t[14] = 44337347
          "10101000100110011001111110" when "00001111", -- t[15] = 44197502
          "10101000000100100100001101" when "00010000", -- t[16] = 44058893
          "10100111100011000001010111" when "00010001", -- t[17] = 43921495
          "10100111000001110001010001" when "00010010", -- t[18] = 43785297
          "10100110100000110011100001" when "00010011", -- t[19] = 43650273
          "10100110000000000111111110" when "00010100", -- t[20] = 43516414
          "10100101011111101110001111" when "00010101", -- t[21] = 43383695
          "10100100111111100110001011" when "00010110", -- t[22] = 43252107
          "10100100011111101111011010" when "00010111", -- t[23] = 43121626
          "10100100000000001001110011" when "00011000", -- t[24] = 42992243
          "10100011100000110100111111" when "00011001", -- t[25] = 42863935
          "10100011000001110000110111" when "00011010", -- t[26] = 42736695
          "10100010100010111101000100" when "00011011", -- t[27] = 42610500
          "10100010000100011001011110" when "00011100", -- t[28] = 42485342
          "10100001100110000101110000" when "00011101", -- t[29] = 42361200
          "10100001001000000001110011" when "00011110", -- t[30] = 42238067
          "10100000101010001101010010" when "00011111", -- t[31] = 42115922
          "10100000001100101000000101" when "00100000", -- t[32] = 41994757
          "10011111101111010001111010" when "00100001", -- t[33] = 41874554
          "10011111010010001010101001" when "00100010", -- t[34] = 41755305
          "10011110110101010010000000" when "00100011", -- t[35] = 41636992
          "10011110011000100111110111" when "00100100", -- t[36] = 41519607
          "10011101111100001011111101" when "00100101", -- t[37] = 41403133
          "10011101011111111110001011" when "00100110", -- t[38] = 41287563
          "10011101000011111110010000" when "00100111", -- t[39] = 41172880
          "10011100101000001100000110" when "00101000", -- t[40] = 41059078
          "10011100001100100111011011" when "00101001", -- t[41] = 40946139
          "10011011110001010000001010" when "00101010", -- t[42] = 40834058
          "10011011010110000110000010" when "00101011", -- t[43] = 40722818
          "10011010111011001000111111" when "00101100", -- t[44] = 40612415
          "10011010100000011000101111" when "00101101", -- t[45] = 40502831
          "10011010000101110101001110" when "00101110", -- t[46] = 40394062
          "10011001101011011110001101" when "00101111", -- t[47] = 40286093
          "10011001010001010011100110" when "00110000", -- t[48] = 40178918
          "10011000110111010101001011" when "00110001", -- t[49] = 40072523
          "10011000011101100010110111" when "00110010", -- t[50] = 39966903
          "10011000000011111100011011" when "00110011", -- t[51] = 39862043
          "10010111101010100001110011" when "00110100", -- t[52] = 39757939
          "10010111010001010010110001" when "00110101", -- t[53] = 39654577
          "10010110111000001111010000" when "00110110", -- t[54] = 39551952
          "10010110011111010111000100" when "00110111", -- t[55] = 39450052
          "10010110000110101010000111" when "00111000", -- t[56] = 39348871
          "10010101101110001000001110" when "00111001", -- t[57] = 39248398
          "10010101010101110001010010" when "00111010", -- t[58] = 39148626
          "10010100111101100101001010" when "00111011", -- t[59] = 39049546
          "10010100100101100011101111" when "00111100", -- t[60] = 38951151
          "10010100001101101100110110" when "00111101", -- t[61] = 38853430
          "10010011110110000000011100" when "00111110", -- t[62] = 38756380
          "10010011011110011110010100" when "00111111", -- t[63] = 38659988
          "10010011000111000110011011" when "01000000", -- t[64] = 38564251
          "10010010101111111000100110" when "01000001", -- t[65] = 38469158
          "10010010011000110100110000" when "01000010", -- t[66] = 38374704
          "10010010000001111010101111" when "01000011", -- t[67] = 38280879
          "10010001101011001010100000" when "01000100", -- t[68] = 38187680
          "10010001010100100011110111" when "01000101", -- t[69] = 38095095
          "10010000111110000110110010" when "01000110", -- t[70] = 38003122
          "10010000100111110011000110" when "01000111", -- t[71] = 37911750
          "10010000010001101000110000" when "01001000", -- t[72] = 37820976
          "10001111111011100111100101" when "01001001", -- t[73] = 37730789
          "10001111100101101111100100" when "01001010", -- t[74] = 37641188
          "10001111010000000000100001" when "01001011", -- t[75] = 37552161
          "10001110111010011010011010" when "01001100", -- t[76] = 37463706
          "10001110100100111101000111" when "01001101", -- t[77] = 37375815
          "10001110001111101000100010" when "01001110", -- t[78] = 37288482
          "10001101111010011100100101" when "01001111", -- t[79] = 37201701
          "10001101100101011001001011" when "01010000", -- t[80] = 37115467
          "10001101010000011110001100" when "01010001", -- t[81] = 37029772
          "10001100111011101011100101" when "01010010", -- t[82] = 36944613
          "10001100100111000001001110" when "01010011", -- t[83] = 36859982
          "10001100010010011111000011" when "01010100", -- t[84] = 36775875
          "10001011111110000100111110" when "01010101", -- t[85] = 36692286
          "10001011101001110010111010" when "01010110", -- t[86] = 36609210
          "10001011010101101000110000" when "01010111", -- t[87] = 36526640
          "10001011000001100110011110" when "01011000", -- t[88] = 36444574
          "10001010101101101011111011" when "01011001", -- t[89] = 36363003
          "10001010011001111001000101" when "01011010", -- t[90] = 36281925
          "10001010000110001101110101" when "01011011", -- t[91] = 36201333
          "10001001110010101010001000" when "01011100", -- t[92] = 36121224
          "10001001011111001101110110" when "01011101", -- t[93] = 36041590
          "10001001001011111000111110" when "01011110", -- t[94] = 35962430
          "10001000111000101011011001" when "01011111", -- t[95] = 35883737
          "10001000100101100101000011" when "01100000", -- t[96] = 35805507
          "10001000010010100101110110" when "01100001", -- t[97] = 35727734
          "10000111111111101101110000" when "01100010", -- t[98] = 35650416
          "10000111101100111100101011" when "01100011", -- t[99] = 35573547
          "10000111011010010010100011" when "01100100", -- t[100] = 35497123
          "10000111000111101111010011" when "01100101", -- t[101] = 35421139
          "10000110110101010010110111" when "01100110", -- t[102] = 35345591
          "10000110100010111101001011" when "01100111", -- t[103] = 35270475
          "10000110010000101110001100" when "01101000", -- t[104] = 35195788
          "10000101111110100101110011" when "01101001", -- t[105] = 35121523
          "10000101101100100011111111" when "01101010", -- t[106] = 35047679
          "10000101011010101000101001" when "01101011", -- t[107] = 34974249
          "10000101001000110011110001" when "01101100", -- t[108] = 34901233
          "10000100110111000101001111" when "01101101", -- t[109] = 34828623
          "10000100100101011101000010" when "01101110", -- t[110] = 34756418
          "10000100010011111011000100" when "01101111", -- t[111] = 34684612
          "10000100000010011111010011" when "01110000", -- t[112] = 34613203
          "10000011110001001001101011" when "01110001", -- t[113] = 34542187
          "10000011011111111010001000" when "01110010", -- t[114] = 34471560
          "10000011001110110000100110" when "01110011", -- t[115] = 34401318
          "10000010111101101101000011" when "01110100", -- t[116] = 34331459
          "10000010101100101111011010" when "01110101", -- t[117] = 34261978
          "10000010011011110111101000" when "01110110", -- t[118] = 34192872
          "10000010001011000101101010" when "01110111", -- t[119] = 34124138
          "10000001111010011001011100" when "01111000", -- t[120] = 34055772
          "10000001101001110010111010" when "01111001", -- t[121] = 33987770
          "10000001011001010010000011" when "01111010", -- t[122] = 33920131
          "10000001001000110110110010" when "01111011", -- t[123] = 33852850
          "10000000111000100001000100" when "01111100", -- t[124] = 33785924
          "10000000101000010000110110" when "01111101", -- t[125] = 33719350
          "10000000011000000110000101" when "01111110", -- t[126] = 33653125
          "10000000001000000000101110" when "01111111", -- t[127] = 33587246
          "01111111111000000000101110" when "10000000", -- t[128] = 33521710
          "01111111101000000110000010" when "10000001", -- t[129] = 33456514
          "01111111011000010000100111" when "10000010", -- t[130] = 33391655
          "01111111001000100000011001" when "10000011", -- t[131] = 33327129
          "01111110111000110101010111" when "10000100", -- t[132] = 33262935
          "01111110101001001111011100" when "10000101", -- t[133] = 33199068
          "01111110011001101110101000" when "10000110", -- t[134] = 33135528
          "01111110001010010010110101" when "10000111", -- t[135] = 33072309
          "01111101111010111100000011" when "10001000", -- t[136] = 33009411
          "01111101101011101010001110" when "10001001", -- t[137] = 32946830
          "01111101011100011101010011" when "10001010", -- t[138] = 32884563
          "01111101001101010101010000" when "10001011", -- t[139] = 32822608
          "01111100111110010010000010" when "10001100", -- t[140] = 32760962
          "01111100101111010011100111" when "10001101", -- t[141] = 32699623
          "01111100100000011001111100" when "10001110", -- t[142] = 32638588
          "01111100010001100100111110" when "10001111", -- t[143] = 32577854
          "01111100000010110100101011" when "10010000", -- t[144] = 32517419
          "01111011110100001001000001" when "10010001", -- t[145] = 32457281
          "01111011100101100001111101" when "10010010", -- t[146] = 32397437
          "01111011010110111111011100" when "10010011", -- t[147] = 32337884
          "01111011001000100001011101" when "10010100", -- t[148] = 32278621
          "01111010111010000111111101" when "10010101", -- t[149] = 32219645
          "01111010101011110010111001" when "10010110", -- t[150] = 32160953
          "01111010011101100010010000" when "10010111", -- t[151] = 32102544
          "01111010001111010101111110" when "10011000", -- t[152] = 32044414
          "01111010000001001110000011" when "10011001", -- t[153] = 31986563
          "01111001110011001010011011" when "10011010", -- t[154] = 31928987
          "01111001100101001011000100" when "10011011", -- t[155] = 31871684
          "01111001010111001111111100" when "10011100", -- t[156] = 31814652
          "01111001001001011001000001" when "10011101", -- t[157] = 31757889
          "01111000111011100110010010" when "10011110", -- t[158] = 31701394
          "01111000101101110111101011" when "10011111", -- t[159] = 31645163
          "01111000100000001101001011" when "10100000", -- t[160] = 31589195
          "01111000010010100110101111" when "10100001", -- t[161] = 31533487
          "01111000000101000100010110" when "10100010", -- t[162] = 31478038
          "01110111110111100101111110" when "10100011", -- t[163] = 31422846
          "01110111101010001011100100" when "10100100", -- t[164] = 31367908
          "01110111011100110101000111" when "10100101", -- t[165] = 31313223
          "01110111001111100010100100" when "10100110", -- t[166] = 31258788
          "01110111000010010011111010" when "10100111", -- t[167] = 31204602
          "01110110110101001001001000" when "10101000", -- t[168] = 31150664
          "01110110101000000010001010" when "10101001", -- t[169] = 31096970
          "01110110011010111110111111" when "10101010", -- t[170] = 31043519
          "01110110001101111111100110" when "10101011", -- t[171] = 30990310
          "01110110000001000011111100" when "10101100", -- t[172] = 30937340
          "01110101110100001011111111" when "10101101", -- t[173] = 30884607
          "01110101100111010111101111" when "10101110", -- t[174] = 30832111
          "01110101011010100111001000" when "10101111", -- t[175] = 30779848
          "01110101001101111010001011" when "10110000", -- t[176] = 30727819
          "01110101000001010000110011" when "10110001", -- t[177] = 30676019
          "01110100110100101011000001" when "10110010", -- t[178] = 30624449
          "01110100101000001000110001" when "10110011", -- t[179] = 30573105
          "01110100011011101010000100" when "10110100", -- t[180] = 30521988
          "01110100001111001110110110" when "10110101", -- t[181] = 30471094
          "01110100000010110111000110" when "10110110", -- t[182] = 30420422
          "01110011110110100010110011" when "10110111", -- t[183] = 30369971
          "01110011101010010001111011" when "10111000", -- t[184] = 30319739
          "01110011011110000100011101" when "10111001", -- t[185] = 30269725
          "01110011010001111010010110" when "10111010", -- t[186] = 30219926
          "01110011000101110011100110" when "10111011", -- t[187] = 30170342
          "01110010111001110000001010" when "10111100", -- t[188] = 30120970
          "01110010101101110000000010" when "10111101", -- t[189] = 30071810
          "01110010100001110011001011" when "10111110", -- t[190] = 30022859
          "01110010010101111001100101" when "10111111", -- t[191] = 29974117
          "01110010001010000011001101" when "11000000", -- t[192] = 29925581
          "01110001111110010000000011" when "11000001", -- t[193] = 29877251
          "01110001110010100000000101" when "11000010", -- t[194] = 29829125
          "01110001100110110011010000" when "11000011", -- t[195] = 29781200
          "01110001011011001001100101" when "11000100", -- t[196] = 29733477
          "01110001001111100011000010" when "11000101", -- t[197] = 29685954
          "01110001000011111111100101" when "11000110", -- t[198] = 29638629
          "01110000111000011111001100" when "11000111", -- t[199] = 29591500
          "01110000101101000001110111" when "11001000", -- t[200] = 29544567
          "01110000100001100111100100" when "11001001", -- t[201] = 29497828
          "01110000010110010000010001" when "11001010", -- t[202] = 29451281
          "01110000001010111011111110" when "11001011", -- t[203] = 29404926
          "01101111111111101010101010" when "11001100", -- t[204] = 29358762
          "01101111110100011100010010" when "11001101", -- t[205] = 29312786
          "01101111101001010000110101" when "11001110", -- t[206] = 29266997
          "01101111011110001000010011" when "11001111", -- t[207] = 29221395
          "01101111010011000010101010" when "11010000", -- t[208] = 29175978
          "01101111000111111111111000" when "11010001", -- t[209] = 29130744
          "01101110111100111111111101" when "11010010", -- t[210] = 29085693
          "01101110110010000010110111" when "11010011", -- t[211] = 29040823
          "01101110100111001000100101" when "11010100", -- t[212] = 28996133
          "01101110011100010001000110" when "11010101", -- t[213] = 28951622
          "01101110010001011100011001" when "11010110", -- t[214] = 28907289
          "01101110000110101010011100" when "11010111", -- t[215] = 28863132
          "01101101111011111011001111" when "11011000", -- t[216] = 28819151
          "01101101110001001110101111" when "11011001", -- t[217] = 28775343
          "01101101100110100100111101" when "11011010", -- t[218] = 28731709
          "01101101011011111101110110" when "11011011", -- t[219] = 28688246
          "01101101010001011001011010" when "11011100", -- t[220] = 28644954
          "01101101000110110111100111" when "11011101", -- t[221] = 28601831
          "01101100111100011000011110" when "11011110", -- t[222] = 28558878
          "01101100110001111011111011" when "11011111", -- t[223] = 28516091
          "01101100100111100001111111" when "11100000", -- t[224] = 28473471
          "01101100011101001010101000" when "11100001", -- t[225] = 28431016
          "01101100010010110101110101" when "11100010", -- t[226] = 28388725
          "01101100001000100011100101" when "11100011", -- t[227] = 28346597
          "01101011111110010011111000" when "11100100", -- t[228] = 28304632
          "01101011110100000110101011" when "11100101", -- t[229] = 28262827
          "01101011101001111011111110" when "11100110", -- t[230] = 28221182
          "01101011011111110011110001" when "11100111", -- t[231] = 28179697
          "01101011010101101110000001" when "11101000", -- t[232] = 28138369
          "01101011001011101010101110" when "11101001", -- t[233] = 28097198
          "01101011000001101001110111" when "11101010", -- t[234] = 28056183
          "01101010110111101011011011" when "11101011", -- t[235] = 28015323
          "01101010101101101111011010" when "11101100", -- t[236] = 27974618
          "01101010100011110101110001" when "11101101", -- t[237] = 27934065
          "01101010011001111110100000" when "11101110", -- t[238] = 27893664
          "01101010010000001001100110" when "11101111", -- t[239] = 27853414
          "01101010000110010111000011" when "11110000", -- t[240] = 27813315
          "01101001111100100110110101" when "11110001", -- t[241] = 27773365
          "01101001110010111000111011" when "11110010", -- t[242] = 27733563
          "01101001101001001101010101" when "11110011", -- t[243] = 27693909
          "01101001011111100100000001" when "11110100", -- t[244] = 27654401
          "01101001010101111100111110" when "11110101", -- t[245] = 27615038
          "01101001001100011000001101" when "11110110", -- t[246] = 27575821
          "01101001000010110101101011" when "11110111", -- t[247] = 27536747
          "01101000111001010101011000" when "11111000", -- t[248] = 27497816
          "01101000101111110111010100" when "11111001", -- t[249] = 27459028
          "01101000100110011011011100" when "11111010", -- t[250] = 27420380
          "01101000011101000001110001" when "11111011", -- t[251] = 27381873
          "01101000010011101010010001" when "11111100", -- t[252] = 27343505
          "01101000001010010100111100" when "11111101", -- t[253] = 27305276
          "01101000000001000001110001" when "11111110", -- t[254] = 27267185
          "01100111110111110000101111" when "11111111", -- t[255] = 27229231
          "--------------------------" when others;

  r(25 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 14; mu_1 = 14; lambda_1 = 14.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t1_pow is
  port ( x : in  std_logic_vector(12 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of fp_log_log_22_t1_pow is
  signal pp0 : std_logic_vector(12 downto 0);
  signal r0 : std_logic_vector(12 downto 0);
begin
  pp0(12) <= x(12);

  pp0(11) <= x(11);

  pp0(10) <= x(10);

  pp0(9) <= x(9);

  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(12 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 8; wO_1,1 = 18.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t1_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(17 downto 0) );
end entity;

architecture arch of fp_log_log_22_t1_t1 is
  signal x : std_logic_vector(7 downto 0);
begin
  x <= a;

  with x select
    r <= "100111000101011100" when "00000000", -- t[0] = 160092
         "100110101101001001" when "00000001", -- t[1] = 158537
         "100110010101001111" when "00000010", -- t[2] = 157007
         "100101111101101110" when "00000011", -- t[3] = 155502
         "100101100110100111" when "00000100", -- t[4] = 154023
         "100101001111110111" when "00000101", -- t[5] = 152567
         "100100111001011111" when "00000110", -- t[6] = 151135
         "100100100011011110" when "00000111", -- t[7] = 149726
         "100100001101110100" when "00001000", -- t[8] = 148340
         "100011111000100000" when "00001001", -- t[9] = 146976
         "100011100011100001" when "00001010", -- t[10] = 145633
         "100011001110110111" when "00001011", -- t[11] = 144311
         "100010111010100010" when "00001100", -- t[12] = 143010
         "100010100110100000" when "00001101", -- t[13] = 141728
         "100010010010110011" when "00001110", -- t[14] = 140467
         "100001111111011000" when "00001111", -- t[15] = 139224
         "100001101100010001" when "00010000", -- t[16] = 138001
         "100001011001011100" when "00010001", -- t[17] = 136796
         "100001000110111001" when "00010010", -- t[18] = 135609
         "100000110100100111" when "00010011", -- t[19] = 134439
         "100000100010100111" when "00010100", -- t[20] = 133287
         "100000010000110111" when "00010101", -- t[21] = 132151
         "011111111111011001" when "00010110", -- t[22] = 131033
         "011111101110001010" when "00010111", -- t[23] = 129930
         "011111011101001011" when "00011000", -- t[24] = 128843
         "011111001100011100" when "00011001", -- t[25] = 127772
         "011110111011111100" when "00011010", -- t[26] = 126716
         "011110101011101011" when "00011011", -- t[27] = 125675
         "011110011011101000" when "00011100", -- t[28] = 124648
         "011110001011110100" when "00011101", -- t[29] = 123636
         "011101111100001101" when "00011110", -- t[30] = 122637
         "011101101100110101" when "00011111", -- t[31] = 121653
         "011101011101101010" when "00100000", -- t[32] = 120682
         "011101001110101100" when "00100001", -- t[33] = 119724
         "011100111111111011" when "00100010", -- t[34] = 118779
         "011100110001010111" when "00100011", -- t[35] = 117847
         "011100100011000000" when "00100100", -- t[36] = 116928
         "011100010100110100" when "00100101", -- t[37] = 116020
         "011100000110110101" when "00100110", -- t[38] = 115125
         "011011111001000001" when "00100111", -- t[39] = 114241
         "011011101011011001" when "00101000", -- t[40] = 113369
         "011011011101111100" when "00101001", -- t[41] = 112508
         "011011010000101011" when "00101010", -- t[42] = 111659
         "011011000011100100" when "00101011", -- t[43] = 110820
         "011010110110101000" when "00101100", -- t[44] = 109992
         "011010101001110111" when "00101101", -- t[45] = 109175
         "011010011101010000" when "00101110", -- t[46] = 108368
         "011010010000110011" when "00101111", -- t[47] = 107571
         "011010000100100000" when "00110000", -- t[48] = 106784
         "011001111000010110" when "00110001", -- t[49] = 106006
         "011001101100010111" when "00110010", -- t[50] = 105239
         "011001100000100001" when "00110011", -- t[51] = 104481
         "011001010100110100" when "00110100", -- t[52] = 103732
         "011001001001010000" when "00110101", -- t[53] = 102992
         "011000111101110101" when "00110110", -- t[54] = 102261
         "011000110010100011" when "00110111", -- t[55] = 101539
         "011000100111011010" when "00111000", -- t[56] = 100826
         "011000011100011001" when "00111001", -- t[57] = 100121
         "011000010001100001" when "00111010", -- t[58] = 99425
         "011000000110110001" when "00111011", -- t[59] = 98737
         "010111111100001001" when "00111100", -- t[60] = 98057
         "010111110001101000" when "00111101", -- t[61] = 97384
         "010111100111010000" when "00111110", -- t[62] = 96720
         "010111011100111111" when "00111111", -- t[63] = 96063
         "010111010010110110" when "01000000", -- t[64] = 95414
         "010111001000110101" when "01000001", -- t[65] = 94773
         "010110111110111010" when "01000010", -- t[66] = 94138
         "010110110101000111" when "01000011", -- t[67] = 93511
         "010110101011011011" when "01000100", -- t[68] = 92891
         "010110100001110110" when "01000101", -- t[69] = 92278
         "010110011000011000" when "01000110", -- t[70] = 91672
         "010110001111000000" when "01000111", -- t[71] = 91072
         "010110000101101111" when "01001000", -- t[72] = 90479
         "010101111100100101" when "01001001", -- t[73] = 89893
         "010101110011100001" when "01001010", -- t[74] = 89313
         "010101101010100100" when "01001011", -- t[75] = 88740
         "010101100001101100" when "01001100", -- t[76] = 88172
         "010101011000111011" when "01001101", -- t[77] = 87611
         "010101010000010000" when "01001110", -- t[78] = 87056
         "010101000111101011" when "01001111", -- t[79] = 86507
         "010100111111001100" when "01010000", -- t[80] = 85964
         "010100110110110010" when "01010001", -- t[81] = 85426
         "010100101110011110" when "01010010", -- t[82] = 84894
         "010100100110010000" when "01010011", -- t[83] = 84368
         "010100011110000111" when "01010100", -- t[84] = 83847
         "010100010110000100" when "01010101", -- t[85] = 83332
         "010100001110000110" when "01010110", -- t[86] = 82822
         "010100000110001101" when "01010111", -- t[87] = 82317
         "010011111110011010" when "01011000", -- t[88] = 81818
         "010011110110101100" when "01011001", -- t[89] = 81324
         "010011101111000010" when "01011010", -- t[90] = 80834
         "010011100111011110" when "01011011", -- t[91] = 80350
         "010011011111111111" when "01011100", -- t[92] = 79871
         "010011011000100100" when "01011101", -- t[93] = 79396
         "010011010001001110" when "01011110", -- t[94] = 78926
         "010011001001111101" when "01011111", -- t[95] = 78461
         "010011000010110001" when "01100000", -- t[96] = 78001
         "010010111011101001" when "01100001", -- t[97] = 77545
         "010010110100100101" when "01100010", -- t[98] = 77093
         "010010101101100110" when "01100011", -- t[99] = 76646
         "010010100110101100" when "01100100", -- t[100] = 76204
         "010010011111110101" when "01100101", -- t[101] = 75765
         "010010011001000011" when "01100110", -- t[102] = 75331
         "010010010010010101" when "01100111", -- t[103] = 74901
         "010010001011101100" when "01101000", -- t[104] = 74476
         "010010000101000110" when "01101001", -- t[105] = 74054
         "010001111110100100" when "01101010", -- t[106] = 73636
         "010001111000000111" when "01101011", -- t[107] = 73223
         "010001110001101101" when "01101100", -- t[108] = 72813
         "010001101011010111" when "01101101", -- t[109] = 72407
         "010001100101000101" when "01101110", -- t[110] = 72005
         "010001011110110111" when "01101111", -- t[111] = 71607
         "010001011000101100" when "01110000", -- t[112] = 71212
         "010001010010100101" when "01110001", -- t[113] = 70821
         "010001001100100010" when "01110010", -- t[114] = 70434
         "010001000110100010" when "01110011", -- t[115] = 70050
         "010001000000100110" when "01110100", -- t[116] = 69670
         "010000111010101101" when "01110101", -- t[117] = 69293
         "010000110100111000" when "01110110", -- t[118] = 68920
         "010000101111000110" when "01110111", -- t[119] = 68550
         "010000101001010111" when "01111000", -- t[120] = 68183
         "010000100011101100" when "01111001", -- t[121] = 67820
         "010000011110000100" when "01111010", -- t[122] = 67460
         "010000011000011111" when "01111011", -- t[123] = 67103
         "010000010010111101" when "01111100", -- t[124] = 66749
         "010000001101011111" when "01111101", -- t[125] = 66399
         "010000001000000100" when "01111110", -- t[126] = 66052
         "010000000010101011" when "01111111", -- t[127] = 65707
         "001111111101010110" when "10000000", -- t[128] = 65366
         "001111111000000011" when "10000001", -- t[129] = 65027
         "001111110010110100" when "10000010", -- t[130] = 64692
         "001111101101101000" when "10000011", -- t[131] = 64360
         "001111101000011110" when "10000100", -- t[132] = 64030
         "001111100011010111" when "10000101", -- t[133] = 63703
         "001111011110010011" when "10000110", -- t[134] = 63379
         "001111011001010010" when "10000111", -- t[135] = 63058
         "001111010100010011" when "10001000", -- t[136] = 62739
         "001111001111011000" when "10001001", -- t[137] = 62424
         "001111001010011111" when "10001010", -- t[138] = 62111
         "001111000101101000" when "10001011", -- t[139] = 61800
         "001111000000110100" when "10001100", -- t[140] = 61492
         "001110111100000011" when "10001101", -- t[141] = 61187
         "001110110111010100" when "10001110", -- t[142] = 60884
         "001110110010101000" when "10001111", -- t[143] = 60584
         "001110101101111110" when "10010000", -- t[144] = 60286
         "001110101001010111" when "10010001", -- t[145] = 59991
         "001110100100110010" when "10010010", -- t[146] = 59698
         "001110100000010000" when "10010011", -- t[147] = 59408
         "001110011011101111" when "10010100", -- t[148] = 59119
         "001110010111010010" when "10010101", -- t[149] = 58834
         "001110010010110110" when "10010110", -- t[150] = 58550
         "001110001110011101" when "10010111", -- t[151] = 58269
         "001110001010000110" when "10011000", -- t[152] = 57990
         "001110000101110010" when "10011001", -- t[153] = 57714
         "001110000001011111" when "10011010", -- t[154] = 57439
         "001101111101001111" when "10011011", -- t[155] = 57167
         "001101111001000001" when "10011100", -- t[156] = 56897
         "001101110100110101" when "10011101", -- t[157] = 56629
         "001101110000101011" when "10011110", -- t[158] = 56363
         "001101101100100011" when "10011111", -- t[159] = 56099
         "001101101000011110" when "10100000", -- t[160] = 55838
         "001101100100011010" when "10100001", -- t[161] = 55578
         "001101100000011000" when "10100010", -- t[162] = 55320
         "001101011100011001" when "10100011", -- t[163] = 55065
         "001101011000011011" when "10100100", -- t[164] = 54811
         "001101010100100000" when "10100101", -- t[165] = 54560
         "001101010000100110" when "10100110", -- t[166] = 54310
         "001101001100101110" when "10100111", -- t[167] = 54062
         "001101001000111000" when "10101000", -- t[168] = 53816
         "001101000101000100" when "10101001", -- t[169] = 53572
         "001101000001010010" when "10101010", -- t[170] = 53330
         "001100111101100001" when "10101011", -- t[171] = 53089
         "001100111001110011" when "10101100", -- t[172] = 52851
         "001100110110000110" when "10101101", -- t[173] = 52614
         "001100110010011011" when "10101110", -- t[174] = 52379
         "001100101110110010" when "10101111", -- t[175] = 52146
         "001100101011001010" when "10110000", -- t[176] = 51914
         "001100100111100101" when "10110001", -- t[177] = 51685
         "001100100100000001" when "10110010", -- t[178] = 51457
         "001100100000011110" when "10110011", -- t[179] = 51230
         "001100011100111110" when "10110100", -- t[180] = 51006
         "001100011001011110" when "10110101", -- t[181] = 50782
         "001100010110000001" when "10110110", -- t[182] = 50561
         "001100010010100101" when "10110111", -- t[183] = 50341
         "001100001111001011" when "10111000", -- t[184] = 50123
         "001100001011110010" when "10111001", -- t[185] = 49906
         "001100001000011011" when "10111010", -- t[186] = 49691
         "001100000101000110" when "10111011", -- t[187] = 49478
         "001100000001110010" when "10111100", -- t[188] = 49266
         "001011111110011111" when "10111101", -- t[189] = 49055
         "001011111011001110" when "10111110", -- t[190] = 48846
         "001011110111111111" when "10111111", -- t[191] = 48639
         "001011110100110001" when "11000000", -- t[192] = 48433
         "001011110001100100" when "11000001", -- t[193] = 48228
         "001011101110011001" when "11000010", -- t[194] = 48025
         "001011101011001111" when "11000011", -- t[195] = 47823
         "001011101000000111" when "11000100", -- t[196] = 47623
         "001011100101000000" when "11000101", -- t[197] = 47424
         "001011100001111011" when "11000110", -- t[198] = 47227
         "001011011110110111" when "11000111", -- t[199] = 47031
         "001011011011110100" when "11001000", -- t[200] = 46836
         "001011011000110011" when "11001001", -- t[201] = 46643
         "001011010101110010" when "11001010", -- t[202] = 46450
         "001011010010110100" when "11001011", -- t[203] = 46260
         "001011001111110110" when "11001100", -- t[204] = 46070
         "001011001100111010" when "11001101", -- t[205] = 45882
         "001011001001111111" when "11001110", -- t[206] = 45695
         "001011000111000110" when "11001111", -- t[207] = 45510
         "001011000100001101" when "11010000", -- t[208] = 45325
         "001011000001010110" when "11010001", -- t[209] = 45142
         "001010111110100000" when "11010010", -- t[210] = 44960
         "001010111011101100" when "11010011", -- t[211] = 44780
         "001010111000111000" when "11010100", -- t[212] = 44600
         "001010110110000110" when "11010101", -- t[213] = 44422
         "001010110011010101" when "11010110", -- t[214] = 44245
         "001010110000100101" when "11010111", -- t[215] = 44069
         "001010101101110110" when "11011000", -- t[216] = 43894
         "001010101011001001" when "11011001", -- t[217] = 43721
         "001010101000011100" when "11011010", -- t[218] = 43548
         "001010100101110001" when "11011011", -- t[219] = 43377
         "001010100011000111" when "11011100", -- t[220] = 43207
         "001010100000011110" when "11011101", -- t[221] = 43038
         "001010011101110110" when "11011110", -- t[222] = 42870
         "001010011011001111" when "11011111", -- t[223] = 42703
         "001010011000101001" when "11100000", -- t[224] = 42537
         "001010010110000101" when "11100001", -- t[225] = 42373
         "001010010011100001" when "11100010", -- t[226] = 42209
         "001010010000111111" when "11100011", -- t[227] = 42047
         "001010001110011101" when "11100100", -- t[228] = 41885
         "001010001011111101" when "11100101", -- t[229] = 41725
         "001010001001011101" when "11100110", -- t[230] = 41565
         "001010000110111111" when "11100111", -- t[231] = 41407
         "001010000100100001" when "11101000", -- t[232] = 41249
         "001010000010000101" when "11101001", -- t[233] = 41093
         "001001111111101001" when "11101010", -- t[234] = 40937
         "001001111101001111" when "11101011", -- t[235] = 40783
         "001001111010110101" when "11101100", -- t[236] = 40629
         "001001111000011101" when "11101101", -- t[237] = 40477
         "001001110110000101" when "11101110", -- t[238] = 40325
         "001001110011101110" when "11101111", -- t[239] = 40174
         "001001110001011001" when "11110000", -- t[240] = 40025
         "001001101111000100" when "11110001", -- t[241] = 39876
         "001001101100110000" when "11110010", -- t[242] = 39728
         "001001101010011101" when "11110011", -- t[243] = 39581
         "001001101000001011" when "11110100", -- t[244] = 39435
         "001001100101111010" when "11110101", -- t[245] = 39290
         "001001100011101010" when "11110110", -- t[246] = 39146
         "001001100001011010" when "11110111", -- t[247] = 39002
         "001001011111001100" when "11111000", -- t[248] = 38860
         "001001011100111110" when "11111001", -- t[249] = 38718
         "001001011010110001" when "11111010", -- t[250] = 38577
         "001001011000100101" when "11111011", -- t[251] = 38437
         "001001010110011010" when "11111100", -- t[252] = 38298
         "001001010100010000" when "11111101", -- t[253] = 38160
         "001001010010000110" when "11111110", -- t[254] = 38022
         "001001001111111110" when "11111111", -- t[255] = 37886
         "------------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 8; beta_1 = 14; lambda_1 = 14;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 8; rho_1,1 = 0; sigma_1,1 = 14; wO_1,1 = 18.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         b : in  std_logic_vector(13 downto 0);
         r : out std_logic_vector(25 downto 0) );
end entity;

architecture arch of fp_log_log_22_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(12 downto 0);
  signal s      : std_logic_vector(13 downto 0);
  component fp_log_log_22_t1_pow is
    port ( x : in  std_logic_vector(12 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  signal a_1    : std_logic_vector(7 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(12 downto 0);
  signal k_1    : std_logic_vector(17 downto 0);
  signal r0_1   : std_logic_vector(32 downto 0);
  signal r_1    : std_logic_vector(25 downto 0);
  component fp_log_log_22_t1_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(17 downto 0) );
  end component;
begin
  sign <= not b(13);
  b0 <= b(12 downto 0) xor (12 downto 0 => sign);

  pow : fp_log_log_22_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(7 downto 0);
  sign_1 <= not s(13);
  s_1 <= s(12 downto 0) xor (12 downto 0 => sign_1);
  t_1 : fp_log_log_22_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(17 downto 0) <=
    r0_1(32 downto 15) xor (32 downto 15 => (not (sign xor sign_1)));
  r_1(25 downto 18) <= (25 downto 18 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 8; mu_2 = 16; lambda_2 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t2_pow is
  port ( x : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_22_t2_pow is
  signal pp0 : std_logic_vector(14 downto 0);
  signal pp1 : std_logic_vector(14 downto 0);
  signal pp2 : std_logic_vector(14 downto 0);
  signal pp3 : std_logic_vector(14 downto 0);
  signal pp4 : std_logic_vector(14 downto 0);
  signal r0 : std_logic_vector(14 downto 0);
begin
  pp0(14) <= '0';
  pp1(14) <= '0';
  pp2(14) <= '0';
  pp3(14) <= '0';
  pp4(14) <= '0';

  pp0(13) <= x(5) and x(6);
  pp1(13) <= x(6);
  pp2(13) <= '0';
  pp3(13) <= '0';
  pp4(13) <= '0';

  pp0(12) <= x(4) and x(6);
  pp1(12) <= '0';
  pp2(12) <= '0';
  pp3(12) <= '0';
  pp4(12) <= '0';

  pp0(11) <= x(3) and x(6);
  pp1(11) <= x(4) and x(5);
  pp2(11) <= x(5);
  pp3(11) <= '0';
  pp4(11) <= '0';

  pp0(10) <= x(2) and x(6);
  pp1(10) <= x(3) and x(5);
  pp2(10) <= '0';
  pp3(10) <= '0';
  pp4(10) <= '0';

  pp0(9) <= x(1) and x(6);
  pp1(9) <= x(2) and x(5);
  pp2(9) <= x(3) and x(4);
  pp3(9) <= x(4);
  pp4(9) <= '0';

  pp0(8) <= x(0) and x(6);
  pp1(8) <= x(1) and x(5);
  pp2(8) <= x(2) and x(4);
  pp3(8) <= '0';
  pp4(8) <= '0';

  pp0(7) <= x(0) and x(5);
  pp1(7) <= x(1) and x(4);
  pp2(7) <= x(2) and x(3);
  pp3(7) <= x(3);
  pp4(7) <= x(6);

  pp0(6) <= x(0) and x(4);
  pp1(6) <= x(1) and x(3);
  pp2(6) <= x(5);
  pp3(6) <= '0';
  pp4(6) <= '0';

  pp0(5) <= x(0) and x(3);
  pp1(5) <= x(1) and x(2);
  pp2(5) <= x(2);
  pp3(5) <= x(4);
  pp4(5) <= '0';

  pp0(4) <= x(0) and x(2);
  pp1(4) <= x(3);
  pp2(4) <= '0';
  pp3(4) <= '0';
  pp4(4) <= '0';

  pp0(3) <= x(0) and x(1);
  pp1(3) <= x(1);
  pp2(3) <= x(2);
  pp3(3) <= '0';
  pp4(3) <= '0';

  pp0(2) <= x(0);
  pp1(2) <= x(1);
  pp2(2) <= '0';
  pp3(2) <= '0';
  pp4(2) <= '0';

  pp0(1) <= '0';
  pp1(1) <= '0';
  pp2(1) <= '0';
  pp3(1) <= '0';
  pp4(1) <= '0';

  pp0(0) <= '0';
  pp1(0) <= '0';
  pp2(0) <= '0';
  pp3(0) <= '0';
  pp4(0) <= '0';

  r0 <= pp0 + pp1 + pp2 + pp3 + pp4;
  r <= "1" & r0(14 downto 4);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 7; wO_2,1 = 9.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t2_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of fp_log_log_22_t2_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "110000101" when "0000000", -- t[0] = 389
         "101111000" when "0000001", -- t[1] = 376
         "101101100" when "0000010", -- t[2] = 364
         "101100000" when "0000011", -- t[3] = 352
         "101010101" when "0000100", -- t[4] = 341
         "101001010" when "0000101", -- t[5] = 330
         "101000000" when "0000110", -- t[6] = 320
         "100110111" when "0000111", -- t[7] = 311
         "100101101" when "0001000", -- t[8] = 301
         "100100100" when "0001001", -- t[9] = 292
         "100011100" when "0001010", -- t[10] = 284
         "100010100" when "0001011", -- t[11] = 276
         "100001100" when "0001100", -- t[12] = 268
         "100000100" when "0001101", -- t[13] = 260
         "011111101" when "0001110", -- t[14] = 253
         "011110110" when "0001111", -- t[15] = 246
         "011101111" when "0010000", -- t[16] = 239
         "011101001" when "0010001", -- t[17] = 233
         "011100011" when "0010010", -- t[18] = 227
         "011011101" when "0010011", -- t[19] = 221
         "011010111" when "0010100", -- t[20] = 215
         "011010010" when "0010101", -- t[21] = 210
         "011001100" when "0010110", -- t[22] = 204
         "011000111" when "0010111", -- t[23] = 199
         "011000010" when "0011000", -- t[24] = 194
         "010111110" when "0011001", -- t[25] = 190
         "010111001" when "0011010", -- t[26] = 185
         "010110100" when "0011011", -- t[27] = 180
         "010110000" when "0011100", -- t[28] = 176
         "010101100" when "0011101", -- t[29] = 172
         "010101000" when "0011110", -- t[30] = 168
         "010100100" when "0011111", -- t[31] = 164
         "010100000" when "0100000", -- t[32] = 160
         "010011101" when "0100001", -- t[33] = 157
         "010011001" when "0100010", -- t[34] = 153
         "010010110" when "0100011", -- t[35] = 150
         "010010011" when "0100100", -- t[36] = 147
         "010001111" when "0100101", -- t[37] = 143
         "010001100" when "0100110", -- t[38] = 140
         "010001001" when "0100111", -- t[39] = 137
         "010000110" when "0101000", -- t[40] = 134
         "010000100" when "0101001", -- t[41] = 132
         "010000001" when "0101010", -- t[42] = 129
         "001111110" when "0101011", -- t[43] = 126
         "001111100" when "0101100", -- t[44] = 124
         "001111001" when "0101101", -- t[45] = 121
         "001110111" when "0101110", -- t[46] = 119
         "001110100" when "0101111", -- t[47] = 116
         "001110010" when "0110000", -- t[48] = 114
         "001110000" when "0110001", -- t[49] = 112
         "001101110" when "0110010", -- t[50] = 110
         "001101011" when "0110011", -- t[51] = 107
         "001101001" when "0110100", -- t[52] = 105
         "001100111" when "0110101", -- t[53] = 103
         "001100101" when "0110110", -- t[54] = 101
         "001100100" when "0110111", -- t[55] = 100
         "001100010" when "0111000", -- t[56] = 98
         "001100000" when "0111001", -- t[57] = 96
         "001011110" when "0111010", -- t[58] = 94
         "001011100" when "0111011", -- t[59] = 92
         "001011011" when "0111100", -- t[60] = 91
         "001011001" when "0111101", -- t[61] = 89
         "001011000" when "0111110", -- t[62] = 88
         "001010110" when "0111111", -- t[63] = 86
         "001010101" when "1000000", -- t[64] = 85
         "001010011" when "1000001", -- t[65] = 83
         "001010010" when "1000010", -- t[66] = 82
         "001010000" when "1000011", -- t[67] = 80
         "001001111" when "1000100", -- t[68] = 79
         "001001110" when "1000101", -- t[69] = 78
         "001001100" when "1000110", -- t[70] = 76
         "001001011" when "1000111", -- t[71] = 75
         "001001010" when "1001000", -- t[72] = 74
         "001001001" when "1001001", -- t[73] = 73
         "001000111" when "1001010", -- t[74] = 71
         "001000110" when "1001011", -- t[75] = 70
         "001000101" when "1001100", -- t[76] = 69
         "001000100" when "1001101", -- t[77] = 68
         "001000011" when "1001110", -- t[78] = 67
         "001000010" when "1001111", -- t[79] = 66
         "001000001" when "1010000", -- t[80] = 65
         "001000000" when "1010001", -- t[81] = 64
         "000111111" when "1010010", -- t[82] = 63
         "000111110" when "1010011", -- t[83] = 62
         "000111101" when "1010100", -- t[84] = 61
         "000111100" when "1010101", -- t[85] = 60
         "000111011" when "1010110", -- t[86] = 59
         "000111010" when "1010111", -- t[87] = 58
         "000111001" when "1011000", -- t[88] = 57
         "000111001" when "1011001", -- t[89] = 57
         "000111000" when "1011010", -- t[90] = 56
         "000110111" when "1011011", -- t[91] = 55
         "000110110" when "1011100", -- t[92] = 54
         "000110101" when "1011101", -- t[93] = 53
         "000110101" when "1011110", -- t[94] = 53
         "000110100" when "1011111", -- t[95] = 52
         "000110011" when "1100000", -- t[96] = 51
         "000110010" when "1100001", -- t[97] = 50
         "000110010" when "1100010", -- t[98] = 50
         "000110001" when "1100011", -- t[99] = 49
         "000110000" when "1100100", -- t[100] = 48
         "000110000" when "1100101", -- t[101] = 48
         "000101111" when "1100110", -- t[102] = 47
         "000101110" when "1100111", -- t[103] = 46
         "000101110" when "1101000", -- t[104] = 46
         "000101101" when "1101001", -- t[105] = 45
         "000101101" when "1101010", -- t[106] = 45
         "000101100" when "1101011", -- t[107] = 44
         "000101011" when "1101100", -- t[108] = 43
         "000101011" when "1101101", -- t[109] = 43
         "000101010" when "1101110", -- t[110] = 42
         "000101010" when "1101111", -- t[111] = 42
         "000101001" when "1110000", -- t[112] = 41
         "000101001" when "1110001", -- t[113] = 41
         "000101000" when "1110010", -- t[114] = 40
         "000101000" when "1110011", -- t[115] = 40
         "000100111" when "1110100", -- t[116] = 39
         "000100111" when "1110101", -- t[117] = 39
         "000100110" when "1110110", -- t[118] = 38
         "000100110" when "1110111", -- t[119] = 38
         "000100101" when "1111000", -- t[120] = 37
         "000100101" when "1111001", -- t[121] = 37
         "000100100" when "1111010", -- t[122] = 36
         "000100100" when "1111011", -- t[123] = 36
         "000100011" when "1111100", -- t[124] = 35
         "000100011" when "1111101", -- t[125] = 35
         "000100011" when "1111110", -- t[126] = 35
         "000100010" when "1111111", -- t[127] = 34
         "---------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_2.
-- Decomposition:
--   alpha_2,2 = 3; sigma'_2,2 = 3; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t2_t2 is
  port ( a : in  std_logic_vector(2 downto 0);
         s : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of fp_log_log_22_t2_t2 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a & s;

  with x select
    r <= "0" when "000000", -- t[0] = 0
         "0" when "000001", -- t[1] = 0
         "0" when "000010", -- t[2] = 0
         "0" when "000011", -- t[3] = 0
         "0" when "000100", -- t[4] = 0
         "0" when "000101", -- t[5] = 0
         "0" when "000110", -- t[6] = 0
         "0" when "000111", -- t[7] = 0
         "0" when "001000", -- t[8] = 0
         "0" when "001001", -- t[9] = 0
         "0" when "001010", -- t[10] = 0
         "0" when "001011", -- t[11] = 0
         "0" when "001100", -- t[12] = 0
         "0" when "001101", -- t[13] = 0
         "0" when "001110", -- t[14] = 0
         "0" when "001111", -- t[15] = 0
         "0" when "010000", -- t[16] = 0
         "0" when "010001", -- t[17] = 0
         "0" when "010010", -- t[18] = 0
         "0" when "010011", -- t[19] = 0
         "0" when "010100", -- t[20] = 0
         "0" when "010101", -- t[21] = 0
         "0" when "010110", -- t[22] = 0
         "0" when "010111", -- t[23] = 0
         "0" when "011000", -- t[24] = 0
         "0" when "011001", -- t[25] = 0
         "0" when "011010", -- t[26] = 0
         "0" when "011011", -- t[27] = 0
         "0" when "011100", -- t[28] = 0
         "0" when "011101", -- t[29] = 0
         "0" when "011110", -- t[30] = 0
         "0" when "011111", -- t[31] = 0
         "0" when "100000", -- t[32] = 0
         "0" when "100001", -- t[33] = 0
         "0" when "100010", -- t[34] = 0
         "0" when "100011", -- t[35] = 0
         "0" when "100100", -- t[36] = 0
         "0" when "100101", -- t[37] = 0
         "0" when "100110", -- t[38] = 0
         "0" when "100111", -- t[39] = 0
         "0" when "101000", -- t[40] = 0
         "0" when "101001", -- t[41] = 0
         "0" when "101010", -- t[42] = 0
         "0" when "101011", -- t[43] = 0
         "0" when "101100", -- t[44] = 0
         "0" when "101101", -- t[45] = 0
         "0" when "101110", -- t[46] = 0
         "0" when "101111", -- t[47] = 0
         "0" when "110000", -- t[48] = 0
         "0" when "110001", -- t[49] = 0
         "0" when "110010", -- t[50] = 0
         "0" when "110011", -- t[51] = 0
         "0" when "110100", -- t[52] = 0
         "0" when "110101", -- t[53] = 0
         "0" when "110110", -- t[54] = 0
         "0" when "110111", -- t[55] = 0
         "0" when "111000", -- t[56] = 0
         "0" when "111001", -- t[57] = 0
         "0" when "111010", -- t[58] = 0
         "0" when "111011", -- t[59] = 0
         "0" when "111100", -- t[60] = 0
         "0" when "111101", -- t[61] = 0
         "0" when "111110", -- t[62] = 0
         "0" when "111111", -- t[63] = 0
         "-" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 7; beta_2 = 8; lambda_2 = 12;  m_2 = 2;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 7; rho_2,1 = 0; sigma_2,1 = 8; wO_2,1 = 9;
--   Q_2,2 (ROM):  alpha_2,2 = 3; rho_2,2 = 8; sigma_2,2 = 4; wO_2,2 = 1.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22_t2 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(25 downto 0) );
end entity;

architecture arch of fp_log_log_22_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(6 downto 0);
  signal s      : std_logic_vector(11 downto 0);
  component fp_log_log_22_t2_pow is
    port ( x : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(6 downto 0);
  signal k_1    : std_logic_vector(8 downto 0);
  signal r0_1   : std_logic_vector(17 downto 0);
  signal r_1    : std_logic_vector(25 downto 0);
  component fp_log_log_22_t2_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  signal a_2    : std_logic_vector(2 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(2 downto 0);
  signal r0_2   : std_logic_vector(0 downto 0);
  signal r_2    : std_logic_vector(25 downto 0);
  component fp_log_log_22_t2_t2 is
    port ( a : in  std_logic_vector(2 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;
begin
  sign <= not b(7);
  b0 <= b(6 downto 0) xor (6 downto 0 => sign);

  pow : fp_log_log_22_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(11);
  s_1 <= s(10 downto 4) xor (10 downto 4 => sign_1);
  t_1 : fp_log_log_22_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(8 downto 0) <=
    r0_1(17 downto 9) xor (17 downto 9 => ((sign_1)));
  r_1(25 downto 9) <= (25 downto 9 => ((sign_1)));

  a_2 <= a(6 downto 4);
  sign_2 <= not s(3);
  s_2 <= s(2 downto 0) xor (2 downto 0 => sign_2);
  t_2 : fp_log_log_22_t2_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(0 downto 0) <=
    r0_2 xor (0 downto 0 => ((sign_2)));
  r_2(25 downto 1) <= (25 downto 1 => ((sign_2)));

  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_22 is
  port ( x : in  std_logic_vector(21 downto 0);
         r : out std_logic_vector(25 downto 0) );
end entity;

architecture arch of fp_log_log_22 is
  signal a_0 : std_logic_vector(7 downto 0);
  signal r_0 : std_logic_vector(25 downto 0);
  component fp_log_log_22_t0 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(25 downto 0) );
  end component;

  signal a_1 : std_logic_vector(7 downto 0);
  signal b_1 : std_logic_vector(13 downto 0);
  signal r_1 : std_logic_vector(25 downto 0);
  component fp_log_log_22_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           b : in  std_logic_vector(13 downto 0);
           r : out std_logic_vector(25 downto 0) );
  end component;

  signal a_2 : std_logic_vector(6 downto 0);
  signal b_2 : std_logic_vector(7 downto 0);
  signal r_2 : std_logic_vector(25 downto 0);
  component fp_log_log_22_t2 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(25 downto 0) );
  end component;

begin
  a_0 <= x(21 downto 14);
  t_0 : fp_log_log_22_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(21 downto 14);
  b_1 <= x(13 downto 0);
  t_1 : fp_log_log_22_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(21 downto 15);
  b_2 <= x(13 downto 6);
  t_2 : fp_log_log_22_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 23; wO = 23.
-- Order-2 polynomial approximation.
-- Decomposition:
--   alpha = 8; beta = 15;
--   T_0 (ROM):     alpha_0 = 8; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 8; beta_1 = 15;
--   T_2 (PowMult): alpha_2 = 7; beta_2 = 10.
-- Guard bits: g = 4.
-- Command line: logfp 23 23 2   rom 8 0   pm 8 15  ah 15 15 15  1 0  8 15 0   pm 7 10  ah 10 16 12  1 1  7 8 0  3 4 8


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 8; beta_0 = 0; wO_0 = 28.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t0 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(27 downto 0) );
end entity;

architecture arch of fp_log_log_23_t0 is
  signal x0   : std_logic_vector(7 downto 0);
  signal r0   : std_logic_vector(27 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "1011000100100011101111000101" when "00000000", -- t[0] = 185744325
          "1011000010001000001001111111" when "00000001", -- t[1] = 185107071
          "1010111111101110000101100100" when "00000010", -- t[2] = 184476004
          "1010111101010101011111101101" when "00000011", -- t[3] = 183850989
          "1010111010111110010111010110" when "00000100", -- t[4] = 183231958
          "1010111000101000101010011110" when "00000101", -- t[5] = 182618782
          "1010110110010100011000000011" when "00000110", -- t[6] = 182011395
          "1010110100000001011110001011" when "00000111", -- t[7] = 181409675
          "1010110001101111111011111000" when "00001000", -- t[8] = 180813560
          "1010101111011111101111010100" when "00001001", -- t[9] = 180222932
          "1010101101010000110111100100" when "00001010", -- t[10] = 179637732
          "1010101011000011010010111000" when "00001011", -- t[11] = 179057848
          "1010101000110111000000010111" when "00001100", -- t[12] = 178483223
          "1010100110101011111110010110" when "00001101", -- t[13] = 177913750
          "1010100100100010001011111111" when "00001110", -- t[14] = 177349375
          "1010100010011001100111101100" when "00001111", -- t[15] = 176789996
          "1010100000010010010000101000" when "00010000", -- t[16] = 176235560
          "1010011110001100000101010001" when "00010001", -- t[17] = 175685969
          "1010011100000111000100110110" when "00010010", -- t[18] = 175141174
          "1010011010000011001101111010" when "00010011", -- t[19] = 174601082
          "1010011000000000011111101011" when "00010100", -- t[20] = 174065643
          "1010010101111110111000110010" when "00010101", -- t[21] = 173534770
          "1010010011111110011000011110" when "00010110", -- t[22] = 173008414
          "1010010001111110111101011100" when "00010111", -- t[23] = 172486492
          "1010010000000000100110111110" when "00011000", -- t[24] = 171968958
          "1010001110000011010011110011" when "00011001", -- t[25] = 171455731
          "1010001100000111000011001111" when "00011010", -- t[26] = 170946767
          "1010001010001011110100000101" when "00011011", -- t[27] = 170441989
          "1010001000010001100101101011" when "00011100", -- t[28] = 169941355
          "1010000110011000010110110110" when "00011101", -- t[29] = 169444790
          "1010000100100000000110111111" when "00011110", -- t[30] = 168952255
          "1010000010101000110100111100" when "00011111", -- t[31] = 168463676
          "1010000000110010100000001000" when "00100000", -- t[32] = 167979016
          "1001111110111101000111011101" when "00100001", -- t[33] = 167498205
          "1001111101001000101010011000" when "00100010", -- t[34] = 167021208
          "1001111011010101000111110100" when "00100011", -- t[35] = 166547956
          "1001111001100010011111010000" when "00100100", -- t[36] = 166078416
          "1001110111110000101111101010" when "00100101", -- t[37] = 165612522
          "1001110101111111111000100001" when "00100110", -- t[38] = 165150241
          "1001110100001111111000110110" when "00100111", -- t[39] = 164691510
          "1001110010100000110000001010" when "00101000", -- t[40] = 164236298
          "1001110000110010011101100001" when "00101001", -- t[41] = 163784545
          "1001101111000101000000011011" when "00101010", -- t[42] = 163336219
          "1001101101011000010111111111" when "00101011", -- t[43] = 162891263
          "1001101011101100100011101111" when "00101100", -- t[44] = 162449647
          "1001101010000001100010110010" when "00101101", -- t[45] = 162011314
          "1001101000010111010100101110" when "00101110", -- t[46] = 161576238
          "1001100110101101111000101011" when "00101111", -- t[47] = 161144363
          "1001100101000101001110001110" when "00110000", -- t[48] = 160715662
          "1001100011011101010100100100" when "00110001", -- t[49] = 160290084
          "1001100001110110001011010001" when "00110010", -- t[50] = 159867601
          "1001100000001111110001100011" when "00110011", -- t[51] = 159448163
          "1001011110101010000111000001" when "00110100", -- t[52] = 159031745
          "1001011101000101001010111010" when "00110101", -- t[53] = 158618298
          "1001011011100000111100110110" when "00110110", -- t[54] = 158207798
          "1001011001111101011100000110" when "00110111", -- t[55] = 157800198
          "1001011000011010101000010010" when "00111000", -- t[56] = 157395474
          "1001010110111000100000101100" when "00111001", -- t[57] = 156993580
          "1001010101010111000100111110" when "00111010", -- t[58] = 156594494
          "1001010011110110010100011101" when "00111011", -- t[59] = 156198173
          "1001010010010110001110110000" when "00111100", -- t[60] = 155804592
          "1001010000110110110011010000" when "00111101", -- t[61] = 155413712
          "1001001111011000000001100101" when "00111110", -- t[62] = 155025509
          "1001001101111001111001000111" when "00111111", -- t[63] = 154639943
          "1001001100011100011001100010" when "01000000", -- t[64] = 154256994
          "1001001010111111100010001101" when "01000001", -- t[65] = 153876621
          "1001001001100011010010110101" when "01000010", -- t[66] = 153498805
          "1001001000000111101010110011" when "01000011", -- t[67] = 153123507
          "1001000110101100101001110100" when "01000100", -- t[68] = 152750708
          "1001000101010010001111010011" when "01000101", -- t[69] = 152380371
          "1001000011111000011010111101" when "01000110", -- t[70] = 152012477
          "1001000010011111001100001110" when "01000111", -- t[71] = 151646990
          "1001000001000110100010110100" when "01001000", -- t[72] = 151283892
          "1000111111101110011110001100" when "01001001", -- t[73] = 150923148
          "1000111110010110111110000100" when "01001010", -- t[74] = 150564740
          "1000111101000000000001111011" when "01001011", -- t[75] = 150208635
          "1000111011101001101001011111" when "01001100", -- t[76] = 149854815
          "1000111010010011110100010001" when "01001101", -- t[77] = 149503249
          "1000111000111110100001111111" when "01001110", -- t[78] = 149153919
          "1000110111101001110010001010" when "01001111", -- t[79] = 148806794
          "1000110110010101100100100001" when "01010000", -- t[80] = 148461857
          "1000110101000001111000100110" when "01010001", -- t[81] = 148119078
          "1000110011101110101110001010" when "01010010", -- t[82] = 147778442
          "1000110010011100000100101110" when "01010011", -- t[83] = 147439918
          "1000110001001001111100000011" when "01010100", -- t[84] = 147103491
          "1000101111111000010011101101" when "01010101", -- t[85] = 146769133
          "1000101110100111001011011101" when "01010110", -- t[86] = 146436829
          "1000101101010110100010110111" when "01010111", -- t[87] = 146106551
          "1000101100000110011001101100" when "01011000", -- t[88] = 145778284
          "1000101010110110101111100010" when "01011001", -- t[89] = 145452002
          "1000101001100111100100001010" when "01011010", -- t[90] = 145127690
          "1000101000011000110111001010" when "01011011", -- t[91] = 144805322
          "1000100111001010101000010100" when "01011100", -- t[92] = 144484884
          "1000100101111100110111010000" when "01011101", -- t[93] = 144166352
          "1000100100101111100011101111" when "01011110", -- t[94] = 143849711
          "1000100011100010101101011001" when "01011111", -- t[95] = 143534937
          "1000100010010110010100000010" when "01100000", -- t[96] = 143222018
          "1000100001001010010111010000" when "01100001", -- t[97] = 142910928
          "1000011111111110110110111000" when "01100010", -- t[98] = 142601656
          "1000011110110011110010100010" when "01100011", -- t[99] = 142294178
          "1000011101101001001010000010" when "01100100", -- t[100] = 141988482
          "1000011100011110111101000001" when "01100101", -- t[101] = 141684545
          "1000011011010101001011010100" when "01100110", -- t[102] = 141382356
          "1000011010001011110100100100" when "01100111", -- t[103] = 141081892
          "1000011001000010111000100110" when "01101000", -- t[104] = 140783142
          "1000010111111010010111000011" when "01101001", -- t[105] = 140486083
          "1000010110110010001111110010" when "01101010", -- t[106] = 140190706
          "1000010101101010100010011101" when "01101011", -- t[107] = 139896989
          "1000010100100011001110111001" when "01101100", -- t[108] = 139604921
          "1000010011011100010100110010" when "01101101", -- t[109] = 139314482
          "1000010010010101110011111110" when "01101110", -- t[110] = 139025662
          "1000010001001111101100000111" when "01101111", -- t[111] = 138738439
          "1000010000001001111101000101" when "01110000", -- t[112] = 138452805
          "1000001111000100100110100011" when "01110001", -- t[113] = 138168739
          "1000001101111111101000011000" when "01110010", -- t[114] = 137886232
          "1000001100111011000010010001" when "01110011", -- t[115] = 137605265
          "1000001011110110110100000100" when "01110100", -- t[116] = 137325828
          "1000001010110010111101011111" when "01110101", -- t[117] = 137047903
          "1000001001101111011110011000" when "01110110", -- t[118] = 136771480
          "1000001000101100010110011110" when "01110111", -- t[119] = 136496542
          "1000000111101001100101100110" when "01111000", -- t[120] = 136223078
          "1000000110100111001011100000" when "01111001", -- t[121] = 135951072
          "1000000101100101001000000011" when "01111010", -- t[122] = 135680515
          "1000000100100011011010111110" when "01111011", -- t[123] = 135411390
          "1000000011100010000100000111" when "01111100", -- t[124] = 135143687
          "1000000010100001000011001111" when "01111101", -- t[125] = 134877391
          "1000000001100000011000001101" when "01111110", -- t[126] = 134612493
          "1000000000100000000010110000" when "01111111", -- t[127] = 134348976
          "0111111111100000000010110000" when "10000000", -- t[128] = 134086832
          "0111111110100000010111111110" when "10000001", -- t[129] = 133826046
          "0111111101100001000010010010" when "10000010", -- t[130] = 133566610
          "0111111100100010000001011011" when "10000011", -- t[131] = 133308507
          "0111111011100011010101010010" when "10000100", -- t[132] = 133051730
          "0111111010100100111101101000" when "10000101", -- t[133] = 132796264
          "0111111001100110111010010110" when "10000110", -- t[134] = 132542102
          "0111111000101001001011001100" when "10000111", -- t[135] = 132289228
          "0111110111101011110000000100" when "10001000", -- t[136] = 132037636
          "0111110110101110101000101110" when "10001001", -- t[137] = 131787310
          "0111110101110001110101000100" when "10001010", -- t[138] = 131538244
          "0111110100110101010100110111" when "10001011", -- t[139] = 131290423
          "0111110011111001001000000001" when "10001100", -- t[140] = 131043841
          "0111110010111101001110010011" when "10001101", -- t[141] = 130798483
          "0111110010000001100111100111" when "10001110", -- t[142] = 130554343
          "0111110001000110010011101111" when "10001111", -- t[143] = 130311407
          "0111110000001011010010100101" when "10010000", -- t[144] = 130069669
          "0111101111010000100011111011" when "10010001", -- t[145] = 129829115
          "0111101110010110000111101100" when "10010010", -- t[146] = 129589740
          "0111101101011011111101101001" when "10010011", -- t[147] = 129351529
          "0111101100100010000101101101" when "10010100", -- t[148] = 129114477
          "0111101011101000011111101011" when "10010101", -- t[149] = 128878571
          "0111101010101111001011011101" when "10010110", -- t[150] = 128643805
          "0111101001110110001000110111" when "10010111", -- t[151] = 128410167
          "0111101000111101010111110010" when "10011000", -- t[152] = 128177650
          "0111101000000100111000000010" when "10011001", -- t[153] = 127946242
          "0111100111001100101001100011" when "10011010", -- t[154] = 127715939
          "0111100110010100101100000111" when "10011011", -- t[155] = 127486727
          "0111100101011100111111101001" when "10011100", -- t[156] = 127258601
          "0111100100100101100011111110" when "10011101", -- t[157] = 127031550
          "0111100011101110011001000000" when "10011110", -- t[158] = 126805568
          "0111100010110111011110100011" when "10011111", -- t[159] = 126580643
          "0111100010000000110100100011" when "10100000", -- t[160] = 126356771
          "0111100001001010011010110100" when "10100001", -- t[161] = 126133940
          "0111100000010100010001010001" when "10100010", -- t[162] = 125912145
          "0111011111011110010111101110" when "10100011", -- t[163] = 125691374
          "0111011110101000101110001000" when "10100100", -- t[164] = 125471624
          "0111011101110011010100010011" when "10100101", -- t[165] = 125252883
          "0111011100111110001010001001" when "10100110", -- t[166] = 125035145
          "0111011100001001001111100010" when "10100111", -- t[167] = 124818402
          "0111011011010100100100010111" when "10101000", -- t[168] = 124602647
          "0111011010100000001000011111" when "10101001", -- t[169] = 124387871
          "0111011001101011111011110101" when "10101010", -- t[170] = 124174069
          "0111011000110111111110001111" when "10101011", -- t[171] = 123961231
          "0111011000000100001111100111" when "10101100", -- t[172] = 123749351
          "0111010111010000101111110101" when "10101101", -- t[173] = 123538421
          "0111010110011101011110110100" when "10101110", -- t[174] = 123328436
          "0111010101101010011100011010" when "10101111", -- t[175] = 123119386
          "0111010100110111101000100010" when "10110000", -- t[176] = 122911266
          "0111010100000101000011000100" when "10110001", -- t[177] = 122704068
          "0111010011010010101011111011" when "10110010", -- t[178] = 122497787
          "0111010010100000100010111101" when "10110011", -- t[179] = 122292413
          "0111010001101110101000000111" when "10110100", -- t[180] = 122087943
          "0111010000111100111011001111" when "10110101", -- t[181] = 121884367
          "0111010000001011011100010001" when "10110110", -- t[182] = 121681681
          "0111001111011010001011000101" when "10110111", -- t[183] = 121479877
          "0111001110101001000111100110" when "10111000", -- t[184] = 121278950
          "0111001101111000010001101011" when "10111001", -- t[185] = 121078891
          "0111001101000111101001010001" when "10111010", -- t[186] = 120879697
          "0111001100010111001110010000" when "10111011", -- t[187] = 120681360
          "0111001011100111000000100010" when "10111100", -- t[188] = 120483874
          "0111001010110111000000000000" when "10111101", -- t[189] = 120287232
          "0111001010000111001100100110" when "10111110", -- t[190] = 120091430
          "0111001001010111100110001100" when "10111111", -- t[191] = 119896460
          "0111001000101000001100101110" when "11000000", -- t[192] = 119702318
          "0111000111111001000000000101" when "11000001", -- t[193] = 119508997
          "0111000111001010000000001011" when "11000010", -- t[194] = 119316491
          "0111000110011011001100111010" when "11000011", -- t[195] = 119124794
          "0111000101101100100110001110" when "11000100", -- t[196] = 118933902
          "0111000100111110001100000000" when "11000101", -- t[197] = 118743808
          "0111000100001111111110001011" when "11000110", -- t[198] = 118554507
          "0111000011100001111100101000" when "11000111", -- t[199] = 118365992
          "0111000010110100000111010100" when "11001000", -- t[200] = 118178260
          "0111000010000110011110000111" when "11001001", -- t[201] = 117991303
          "0111000001011001000000111111" when "11001010", -- t[202] = 117805119
          "0111000000101011101111110010" when "11001011", -- t[203] = 117619698
          "0110111111111110101010100000" when "11001100", -- t[204] = 117435040
          "0110111111010001110000111111" when "11001101", -- t[205] = 117251135
          "0110111110100101000011001110" when "11001110", -- t[206] = 117067982
          "0110111101111000100001000100" when "11001111", -- t[207] = 116885572
          "0110111101001100001010100000" when "11010000", -- t[208] = 116703904
          "0110111100011111111111011001" when "11010001", -- t[209] = 116522969
          "0110111011110011111111101101" when "11010010", -- t[210] = 116342765
          "0110111011001000001011010101" when "11010011", -- t[211] = 116163285
          "0110111010011100100010001110" when "11010100", -- t[212] = 115984526
          "0110111001110001000100010010" when "11010101", -- t[213] = 115806482
          "0110111001000101110001011101" when "11010110", -- t[214] = 115629149
          "0110111000011010101001101001" when "11010111", -- t[215] = 115452521
          "0110110111101111101100110011" when "11011000", -- t[216] = 115276595
          "0110110111000100111010110101" when "11011001", -- t[217] = 115101365
          "0110110110011010010011101011" when "11011010", -- t[218] = 114926827
          "0110110101101111110111010000" when "11011011", -- t[219] = 114752976
          "0110110101000101100101100001" when "11011100", -- t[220] = 114579809
          "0110110100011011011110010111" when "11011101", -- t[221] = 114407319
          "0110110011110001100001110000" when "11011110", -- t[222] = 114235504
          "0110110011000111101111100101" when "11011111", -- t[223] = 114064357
          "0110110010011110000111110101" when "11100000", -- t[224] = 113893877
          "0110110001110100101010011001" when "11100001", -- t[225] = 113724057
          "0110110001001011010111001110" when "11100010", -- t[226] = 113554894
          "0110110000100010001110001110" when "11100011", -- t[227] = 113386382
          "0110101111111001001111011000" when "11100100", -- t[228] = 113218520
          "0110101111010000011010100101" when "11100101", -- t[229] = 113051301
          "0110101110100111101111110011" when "11100110", -- t[230] = 112884723
          "0110101101111111001110111100" when "11100111", -- t[231] = 112718780
          "0110101101010110110111111101" when "11101000", -- t[232] = 112553469
          "0110101100101110101010110010" when "11101001", -- t[233] = 112388786
          "0110101100000110100111010111" when "11101010", -- t[234] = 112224727
          "0110101011011110101101100111" when "11101011", -- t[235] = 112061287
          "0110101010110110111101100000" when "11101100", -- t[236] = 111898464
          "0110101010001111010110111100" when "11101101", -- t[237] = 111736252
          "0110101001100111111001111010" when "11101110", -- t[238] = 111574650
          "0110101001000000100110010011" when "11101111", -- t[239] = 111413651
          "0110101000011001011100000110" when "11110000", -- t[240] = 111253254
          "0110100111110010011011001101" when "11110001", -- t[241] = 111093453
          "0110100111001011100011100110" when "11110010", -- t[242] = 110934246
          "0110100110100100110101001100" when "11110011", -- t[243] = 110775628
          "0110100101111110001111111100" when "11110100", -- t[244] = 110617596
          "0110100101010111110011110011" when "11110101", -- t[245] = 110460147
          "0110100100110001100000101101" when "11110110", -- t[246] = 110303277
          "0110100100001011010110100110" when "11110111", -- t[247] = 110146982
          "0110100011100101010101011011" when "11111000", -- t[248] = 109991259
          "0110100010111111011101001000" when "11111001", -- t[249] = 109836104
          "0110100010011001101101101010" when "11111010", -- t[250] = 109681514
          "0110100001110100000110111101" when "11111011", -- t[251] = 109527485
          "0110100001001110101000111111" when "11111100", -- t[252] = 109374015
          "0110100000101001010011101011" when "11111101", -- t[253] = 109221099
          "0110100000000100000110111111" when "11111110", -- t[254] = 109068735
          "0110011111011111000010110110" when "11111111", -- t[255] = 108916918
          "----------------------------" when others;

  r(27 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 15; mu_1 = 15; lambda_1 = 15.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t1_pow is
  port ( x : in  std_logic_vector(13 downto 0);
         r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of fp_log_log_23_t1_pow is
  signal pp0 : std_logic_vector(13 downto 0);
  signal r0 : std_logic_vector(13 downto 0);
begin
  pp0(13) <= x(13);

  pp0(12) <= x(12);

  pp0(11) <= x(11);

  pp0(10) <= x(10);

  pp0(9) <= x(9);

  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(13 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 8; wO_1,1 = 20.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t1_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(19 downto 0) );
end entity;

architecture arch of fp_log_log_23_t1_t1 is
  signal x : std_logic_vector(7 downto 0);
begin
  x <= a;

  with x select
    r <= "10011100010101110001" when "00000000", -- t[0] = 640369
         "10011010110100100010" when "00000001", -- t[1] = 634146
         "10011001010100111011" when "00000010", -- t[2] = 628027
         "10010111110110111010" when "00000011", -- t[3] = 622010
         "10010110011010011011" when "00000100", -- t[4] = 616091
         "10010100111111011101" when "00000101", -- t[5] = 610269
         "10010011100101111101" when "00000110", -- t[6] = 604541
         "10010010001101111001" when "00000111", -- t[7] = 598905
         "10010000110111010000" when "00001000", -- t[8] = 593360
         "10001111100001111110" when "00001001", -- t[9] = 587902
         "10001110001110000011" when "00001010", -- t[10] = 582531
         "10001100111011011011" when "00001011", -- t[11] = 577243
         "10001011101010000110" when "00001100", -- t[12] = 572038
         "10001010011010000001" when "00001101", -- t[13] = 566913
         "10001001001011001011" when "00001110", -- t[14] = 561867
         "10000111111101100010" when "00001111", -- t[15] = 556898
         "10000110110001000011" when "00010000", -- t[16] = 552003
         "10000101100101101111" when "00010001", -- t[17] = 547183
         "10000100011011100010" when "00010010", -- t[18] = 542434
         "10000011010010011100" when "00010011", -- t[19] = 537756
         "10000010001010011011" when "00010100", -- t[20] = 533147
         "10000001000011011110" when "00010101", -- t[21] = 528606
         "01111111111101100010" when "00010110", -- t[22] = 524130
         "01111110111000100111" when "00010111", -- t[23] = 519719
         "01111101110100101100" when "00011000", -- t[24] = 515372
         "01111100110001101111" when "00011001", -- t[25] = 511087
         "01111011101111101111" when "00011010", -- t[26] = 506863
         "01111010101110101010" when "00011011", -- t[27] = 502698
         "01111001101110100000" when "00011100", -- t[28] = 498592
         "01111000101111001111" when "00011101", -- t[29] = 494543
         "01110111110000110110" when "00011110", -- t[30] = 490550
         "01110110110011010100" when "00011111", -- t[31] = 486612
         "01110101110110101000" when "00100000", -- t[32] = 482728
         "01110100111010110001" when "00100001", -- t[33] = 478897
         "01110011111111101110" when "00100010", -- t[34] = 475118
         "01110011000101011101" when "00100011", -- t[35] = 471389
         "01110010001011111111" when "00100100", -- t[36] = 467711
         "01110001010011010001" when "00100101", -- t[37] = 464081
         "01110000011011010011" when "00100110", -- t[38] = 460499
         "01101111100100000101" when "00100111", -- t[39] = 456965
         "01101110101101100101" when "00101000", -- t[40] = 453477
         "01101101110111110010" when "00101001", -- t[41] = 450034
         "01101101000010101011" when "00101010", -- t[42] = 446635
         "01101100001110010000" when "00101011", -- t[43] = 443280
         "01101011011010100000" when "00101100", -- t[44] = 439968
         "01101010100111011011" when "00101101", -- t[45] = 436699
         "01101001110100111110" when "00101110", -- t[46] = 433470
         "01101001000011001010" when "00101111", -- t[47] = 430282
         "01101000010001111110" when "00110000", -- t[48] = 427134
         "01100111100001011010" when "00110001", -- t[49] = 424026
         "01100110110001011011" when "00110010", -- t[50] = 420955
         "01100110000010000011" when "00110011", -- t[51] = 417923
         "01100101010011001111" when "00110100", -- t[52] = 414927
         "01100100100101000000" when "00110101", -- t[53] = 411968
         "01100011110111010101" when "00110110", -- t[54] = 409045
         "01100011001010001110" when "00110111", -- t[55] = 406158
         "01100010011101101000" when "00111000", -- t[56] = 403304
         "01100001110001100101" when "00111001", -- t[57] = 400485
         "01100001000110000011" when "00111010", -- t[58] = 397699
         "01100000011011000011" when "00111011", -- t[59] = 394947
         "01011111110000100010" when "00111100", -- t[60] = 392226
         "01011111000110100001" when "00111101", -- t[61] = 389537
         "01011110011101000000" when "00111110", -- t[62] = 386880
         "01011101110011111101" when "00111111", -- t[63] = 384253
         "01011101001011011001" when "01000000", -- t[64] = 381657
         "01011100100011010010" when "01000001", -- t[65] = 379090
         "01011011111011101001" when "01000010", -- t[66] = 376553
         "01011011010100011100" when "01000011", -- t[67] = 374044
         "01011010101101101100" when "01000100", -- t[68] = 371564
         "01011010000111011000" when "01000101", -- t[69] = 369112
         "01011001100001011111" when "01000110", -- t[70] = 366687
         "01011000111100000001" when "01000111", -- t[71] = 364289
         "01011000010110111110" when "01001000", -- t[72] = 361918
         "01010111110010010100" when "01001001", -- t[73] = 359572
         "01010111001110000101" when "01001010", -- t[74] = 357253
         "01010110101010001111" when "01001011", -- t[75] = 354959
         "01010110000110110010" when "01001100", -- t[76] = 352690
         "01010101100011101101" when "01001101", -- t[77] = 350445
         "01010101000001000000" when "01001110", -- t[78] = 348224
         "01010100011110101100" when "01001111", -- t[79] = 346028
         "01010011111100101111" when "01010000", -- t[80] = 343855
         "01010011011011001001" when "01010001", -- t[81] = 341705
         "01010010111001111001" when "01010010", -- t[82] = 339577
         "01010010011001000000" when "01010011", -- t[83] = 337472
         "01010001111000011101" when "01010100", -- t[84] = 335389
         "01010001011000010000" when "01010101", -- t[85] = 333328
         "01010000111000011000" when "01010110", -- t[86] = 331288
         "01010000011000110110" when "01010111", -- t[87] = 329270
         "01001111111001101000" when "01011000", -- t[88] = 327272
         "01001111011010101110" when "01011001", -- t[89] = 325294
         "01001110111100001001" when "01011010", -- t[90] = 323337
         "01001110011101111000" when "01011011", -- t[91] = 321400
         "01001101111111111010" when "01011100", -- t[92] = 319482
         "01001101100010010000" when "01011101", -- t[93] = 317584
         "01001101000100111001" when "01011110", -- t[94] = 315705
         "01001100100111110100" when "01011111", -- t[95] = 313844
         "01001100001011000010" when "01100000", -- t[96] = 312002
         "01001011101110100010" when "01100001", -- t[97] = 310178
         "01001011010010010101" when "01100010", -- t[98] = 308373
         "01001010110110011001" when "01100011", -- t[99] = 306585
         "01001010011010101110" when "01100100", -- t[100] = 304814
         "01001001111111010101" when "01100101", -- t[101] = 303061
         "01001001100100001101" when "01100110", -- t[102] = 301325
         "01001001001001010101" when "01100111", -- t[103] = 299605
         "01001000101110101110" when "01101000", -- t[104] = 297902
         "01001000010100010111" when "01101001", -- t[105] = 296215
         "01000111111010010001" when "01101010", -- t[106] = 294545
         "01000111100000011010" when "01101011", -- t[107] = 292890
         "01000111000110110011" when "01101100", -- t[108] = 291251
         "01000110101101011100" when "01101101", -- t[109] = 289628
         "01000110010100010100" when "01101110", -- t[110] = 288020
         "01000101111011011010" when "01101111", -- t[111] = 286426
         "01000101100010110000" when "01110000", -- t[112] = 284848
         "01000101001010010100" when "01110001", -- t[113] = 283284
         "01000100110010000111" when "01110010", -- t[114] = 281735
         "01000100011010001000" when "01110011", -- t[115] = 280200
         "01000100000010010111" when "01110100", -- t[116] = 278679
         "01000011101010110100" when "01110101", -- t[117] = 277172
         "01000011010011011111" when "01110110", -- t[118] = 275679
         "01000010111100010111" when "01110111", -- t[119] = 274199
         "01000010100101011101" when "01111000", -- t[120] = 272733
         "01000010001110110000" when "01111001", -- t[121] = 271280
         "01000001111000010000" when "01111010", -- t[122] = 269840
         "01000001100001111100" when "01111011", -- t[123] = 268412
         "01000001001011110110" when "01111100", -- t[124] = 266998
         "01000000110101111100" when "01111101", -- t[125] = 265596
         "01000000100000001110" when "01111110", -- t[126] = 264206
         "01000000001010101101" when "01111111", -- t[127] = 262829
         "00111111110101010111" when "10000000", -- t[128] = 261463
         "00111111100000001110" when "10000001", -- t[129] = 260110
         "00111111001011010000" when "10000010", -- t[130] = 258768
         "00111110110110011110" when "10000011", -- t[131] = 257438
         "00111110100001111000" when "10000100", -- t[132] = 256120
         "00111110001101011100" when "10000101", -- t[133] = 254812
         "00111101111001001101" when "10000110", -- t[134] = 253517
         "00111101100101001000" when "10000111", -- t[135] = 252232
         "00111101010001001110" when "10001000", -- t[136] = 250958
         "00111100111101011111" when "10001001", -- t[137] = 249695
         "00111100101001111010" when "10001010", -- t[138] = 248442
         "00111100010110100000" when "10001011", -- t[139] = 247200
         "00111100000011010001" when "10001100", -- t[140] = 245969
         "00111011110000001100" when "10001101", -- t[141] = 244748
         "00111011011101010001" when "10001110", -- t[142] = 243537
         "00111011001010100000" when "10001111", -- t[143] = 242336
         "00111010110111111001" when "10010000", -- t[144] = 241145
         "00111010100101011011" when "10010001", -- t[145] = 239963
         "00111010010011001000" when "10010010", -- t[146] = 238792
         "00111010000000111110" when "10010011", -- t[147] = 237630
         "00111001101110111110" when "10010100", -- t[148] = 236478
         "00111001011101000111" when "10010101", -- t[149] = 235335
         "00111001001011011001" when "10010110", -- t[150] = 234201
         "00111000111001110100" when "10010111", -- t[151] = 233076
         "00111000101000011001" when "10011000", -- t[152] = 231961
         "00111000010111000110" when "10011001", -- t[153] = 230854
         "00111000000101111101" when "10011010", -- t[154] = 229757
         "00110111110100111100" when "10011011", -- t[155] = 228668
         "00110111100100000011" when "10011100", -- t[156] = 227587
         "00110111010011010100" when "10011101", -- t[157] = 226516
         "00110111000010101100" when "10011110", -- t[158] = 225452
         "00110110110010001101" when "10011111", -- t[159] = 224397
         "00110110100001110111" when "10100000", -- t[160] = 223351
         "00110110010001101000" when "10100001", -- t[161] = 222312
         "00110110000001100010" when "10100010", -- t[162] = 221282
         "00110101110001100011" when "10100011", -- t[163] = 220259
         "00110101100001101101" when "10100100", -- t[164] = 219245
         "00110101010001111110" when "10100101", -- t[165] = 218238
         "00110101000010010111" when "10100110", -- t[166] = 217239
         "00110100110010111000" when "10100111", -- t[167] = 216248
         "00110100100011100000" when "10101000", -- t[168] = 215264
         "00110100010100010000" when "10101001", -- t[169] = 214288
         "00110100000101000111" when "10101010", -- t[170] = 213319
         "00110011110110000110" when "10101011", -- t[171] = 212358
         "00110011100111001100" when "10101100", -- t[172] = 211404
         "00110011011000011001" when "10101101", -- t[173] = 210457
         "00110011001001101101" when "10101110", -- t[174] = 209517
         "00110010111011001000" when "10101111", -- t[175] = 208584
         "00110010101100101010" when "10110000", -- t[176] = 207658
         "00110010011110010011" when "10110001", -- t[177] = 206739
         "00110010010000000011" when "10110010", -- t[178] = 205827
         "00110010000001111001" when "10110011", -- t[179] = 204921
         "00110001110011110110" when "10110100", -- t[180] = 204022
         "00110001100101111010" when "10110101", -- t[181] = 203130
         "00110001011000000100" when "10110110", -- t[182] = 202244
         "00110001001010010101" when "10110111", -- t[183] = 201365
         "00110000111100101100" when "10111000", -- t[184] = 200492
         "00110000101111001001" when "10111001", -- t[185] = 199625
         "00110000100001101101" when "10111010", -- t[186] = 198765
         "00110000010100010111" when "10111011", -- t[187] = 197911
         "00110000000111000111" when "10111100", -- t[188] = 197063
         "00101111111001111101" when "10111101", -- t[189] = 196221
         "00101111101100111001" when "10111110", -- t[190] = 195385
         "00101111011111111011" when "10111111", -- t[191] = 194555
         "00101111010011000011" when "11000000", -- t[192] = 193731
         "00101111000110010001" when "11000001", -- t[193] = 192913
         "00101110111001100100" when "11000010", -- t[194] = 192100
         "00101110101100111110" when "11000011", -- t[195] = 191294
         "00101110100000011101" when "11000100", -- t[196] = 190493
         "00101110010100000001" when "11000101", -- t[197] = 189697
         "00101110000111101011" when "11000110", -- t[198] = 188907
         "00101101111011011011" when "11000111", -- t[199] = 188123
         "00101101101111010000" when "11001000", -- t[200] = 187344
         "00101101100011001010" when "11001001", -- t[201] = 186570
         "00101101010111001010" when "11001010", -- t[202] = 185802
         "00101101001011001111" when "11001011", -- t[203] = 185039
         "00101100111111011001" when "11001100", -- t[204] = 184281
         "00101100110011101000" when "11001101", -- t[205] = 183528
         "00101100100111111101" when "11001110", -- t[206] = 182781
         "00101100011100010110" when "11001111", -- t[207] = 182038
         "00101100010000110101" when "11010000", -- t[208] = 181301
         "00101100000101011001" when "11010001", -- t[209] = 180569
         "00101011111010000001" when "11010010", -- t[210] = 179841
         "00101011101110101111" when "11010011", -- t[211] = 179119
         "00101011100011100001" when "11010100", -- t[212] = 178401
         "00101011011000011000" when "11010101", -- t[213] = 177688
         "00101011001101010100" when "11010110", -- t[214] = 176980
         "00101011000010010100" when "11010111", -- t[215] = 176276
         "00101010110111011010" when "11011000", -- t[216] = 175578
         "00101010101100100011" when "11011001", -- t[217] = 174883
         "00101010100001110010" when "11011010", -- t[218] = 174194
         "00101010010111000101" when "11011011", -- t[219] = 173509
         "00101010001100011100" when "11011100", -- t[220] = 172828
         "00101010000001111000" when "11011101", -- t[221] = 172152
         "00101001110111011000" when "11011110", -- t[222] = 171480
         "00101001101100111101" when "11011111", -- t[223] = 170813
         "00101001100010100110" when "11100000", -- t[224] = 170150
         "00101001011000010011" when "11100001", -- t[225] = 169491
         "00101001001110000100" when "11100010", -- t[226] = 168836
         "00101001000011111010" when "11100011", -- t[227] = 168186
         "00101000111001110100" when "11100100", -- t[228] = 167540
         "00101000101111110010" when "11100101", -- t[229] = 166898
         "00101000100101110100" when "11100110", -- t[230] = 166260
         "00101000011011111010" when "11100111", -- t[231] = 165626
         "00101000010010000101" when "11101000", -- t[232] = 164997
         "00101000001000010011" when "11101001", -- t[233] = 164371
         "00100111111110100101" when "11101010", -- t[234] = 163749
         "00100111110100111011" when "11101011", -- t[235] = 163131
         "00100111101011010101" when "11101100", -- t[236] = 162517
         "00100111100001110011" when "11101101", -- t[237] = 161907
         "00100111011000010100" when "11101110", -- t[238] = 161300
         "00100111001110111010" when "11101111", -- t[239] = 160698
         "00100111000101100011" when "11110000", -- t[240] = 160099
         "00100110111100001111" when "11110001", -- t[241] = 159503
         "00100110110011000000" when "11110010", -- t[242] = 158912
         "00100110101001110100" when "11110011", -- t[243] = 158324
         "00100110100000101100" when "11110100", -- t[244] = 157740
         "00100110010111100111" when "11110101", -- t[245] = 157159
         "00100110001110100110" when "11110110", -- t[246] = 156582
         "00100110000101101001" when "11110111", -- t[247] = 156009
         "00100101111100101111" when "11111000", -- t[248] = 155439
         "00100101110011111000" when "11111001", -- t[249] = 154872
         "00100101101011000101" when "11111010", -- t[250] = 154309
         "00100101100010010101" when "11111011", -- t[251] = 153749
         "00100101011001101001" when "11111100", -- t[252] = 153193
         "00100101010001000000" when "11111101", -- t[253] = 152640
         "00100101001000011010" when "11111110", -- t[254] = 152090
         "00100100111111110111" when "11111111", -- t[255] = 151543
         "--------------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 8; beta_1 = 15; lambda_1 = 15;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 8; rho_1,1 = 0; sigma_1,1 = 15; wO_1,1 = 20.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         b : in  std_logic_vector(14 downto 0);
         r : out std_logic_vector(27 downto 0) );
end entity;

architecture arch of fp_log_log_23_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(13 downto 0);
  signal s      : std_logic_vector(14 downto 0);
  component fp_log_log_23_t1_pow is
    port ( x : in  std_logic_vector(13 downto 0);
           r : out std_logic_vector(14 downto 0) );
  end component;

  signal a_1    : std_logic_vector(7 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(13 downto 0);
  signal k_1    : std_logic_vector(19 downto 0);
  signal r0_1   : std_logic_vector(35 downto 0);
  signal r_1    : std_logic_vector(27 downto 0);
  component fp_log_log_23_t1_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(19 downto 0) );
  end component;
begin
  sign <= not b(14);
  b0 <= b(13 downto 0) xor (13 downto 0 => sign);

  pow : fp_log_log_23_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(7 downto 0);
  sign_1 <= not s(14);
  s_1 <= s(13 downto 0) xor (13 downto 0 => sign_1);
  t_1 : fp_log_log_23_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(19 downto 0) <=
    r0_1(35 downto 16) xor (35 downto 16 => (not (sign xor sign_1)));
  r_1(27 downto 20) <= (27 downto 20 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 10; mu_2 = 16; lambda_2 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t2_pow is
  port ( x : in  std_logic_vector(8 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_23_t2_pow is
  signal pp0 : std_logic_vector(14 downto 0);
  signal pp1 : std_logic_vector(14 downto 0);
  signal pp2 : std_logic_vector(14 downto 0);
  signal pp3 : std_logic_vector(14 downto 0);
  signal pp4 : std_logic_vector(14 downto 0);
  signal pp5 : std_logic_vector(14 downto 0);
  signal r0 : std_logic_vector(14 downto 0);
begin
  pp0(14) <= '0';
  pp1(14) <= '0';
  pp2(14) <= '0';
  pp3(14) <= '0';
  pp4(14) <= '0';
  pp5(14) <= '0';

  pp0(13) <= x(7) and x(8);
  pp1(13) <= x(8);
  pp2(13) <= '0';
  pp3(13) <= '0';
  pp4(13) <= '0';
  pp5(13) <= '0';

  pp0(12) <= x(6) and x(8);
  pp1(12) <= '0';
  pp2(12) <= '0';
  pp3(12) <= '0';
  pp4(12) <= '0';
  pp5(12) <= '0';

  pp0(11) <= x(5) and x(8);
  pp1(11) <= x(6) and x(7);
  pp2(11) <= x(7);
  pp3(11) <= '0';
  pp4(11) <= '0';
  pp5(11) <= '0';

  pp0(10) <= x(4) and x(8);
  pp1(10) <= x(5) and x(7);
  pp2(10) <= '0';
  pp3(10) <= '0';
  pp4(10) <= '0';
  pp5(10) <= '0';

  pp0(9) <= x(3) and x(8);
  pp1(9) <= x(4) and x(7);
  pp2(9) <= x(5) and x(6);
  pp3(9) <= x(6);
  pp4(9) <= '0';
  pp5(9) <= '0';

  pp0(8) <= x(2) and x(8);
  pp1(8) <= x(3) and x(7);
  pp2(8) <= x(4) and x(6);
  pp3(8) <= '0';
  pp4(8) <= '0';
  pp5(8) <= '0';

  pp0(7) <= x(1) and x(8);
  pp1(7) <= x(2) and x(7);
  pp2(7) <= x(3) and x(6);
  pp3(7) <= x(4) and x(5);
  pp4(7) <= x(5);
  pp5(7) <= '0';

  pp0(6) <= x(0) and x(8);
  pp1(6) <= x(1) and x(7);
  pp2(6) <= x(2) and x(6);
  pp3(6) <= x(3) and x(5);
  pp4(6) <= '0';
  pp5(6) <= '0';

  pp0(5) <= x(0) and x(7);
  pp1(5) <= x(1) and x(6);
  pp2(5) <= x(2) and x(5);
  pp3(5) <= x(3) and x(4);
  pp4(5) <= x(4);
  pp5(5) <= x(8);

  pp0(4) <= x(0) and x(6);
  pp1(4) <= x(1) and x(5);
  pp2(4) <= x(2) and x(4);
  pp3(4) <= x(7);
  pp4(4) <= '0';
  pp5(4) <= '0';

  pp0(3) <= x(0) and x(5);
  pp1(3) <= x(1) and x(4);
  pp2(3) <= x(2) and x(3);
  pp3(3) <= x(3);
  pp4(3) <= x(6);
  pp5(3) <= '0';

  pp0(2) <= x(0) and x(4);
  pp1(2) <= x(1) and x(3);
  pp2(2) <= x(5);
  pp3(2) <= '0';
  pp4(2) <= '0';
  pp5(2) <= '0';

  pp0(1) <= x(0) and x(3);
  pp1(1) <= x(1) and x(2);
  pp2(1) <= x(2);
  pp3(1) <= x(4);
  pp4(1) <= '0';
  pp5(1) <= '0';

  pp0(0) <= x(0) and x(2);
  pp1(0) <= x(3);
  pp2(0) <= '0';
  pp3(0) <= '0';
  pp4(0) <= '0';
  pp5(0) <= '0';

  r0 <= pp0 + pp1 + pp2 + pp3 + pp4 + pp5;
  r <= "1" & r0(14 downto 4);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 7; wO_2,1 = 11.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t2_t1 is
  port ( a : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of fp_log_log_23_t2_t1 is
  signal x : std_logic_vector(6 downto 0);
begin
  x <= a;

  with x select
    r <= "11000010100" when "0000000", -- t[0] = 1556
         "10111100000" when "0000001", -- t[1] = 1504
         "10110110000" when "0000010", -- t[2] = 1456
         "10110000001" when "0000011", -- t[3] = 1409
         "10101010100" when "0000100", -- t[4] = 1364
         "10100101010" when "0000101", -- t[5] = 1322
         "10100000001" when "0000110", -- t[6] = 1281
         "10011011010" when "0000111", -- t[7] = 1242
         "10010110101" when "0001000", -- t[8] = 1205
         "10010010010" when "0001001", -- t[9] = 1170
         "10001101111" when "0001010", -- t[10] = 1135
         "10001001111" when "0001011", -- t[11] = 1103
         "10000101111" when "0001100", -- t[12] = 1071
         "10000010001" when "0001101", -- t[13] = 1041
         "01111110100" when "0001110", -- t[14] = 1012
         "01111011000" when "0001111", -- t[15] = 984
         "01110111110" when "0010000", -- t[16] = 958
         "01110100100" when "0010001", -- t[17] = 932
         "01110001011" when "0010010", -- t[18] = 907
         "01101110100" when "0010011", -- t[19] = 884
         "01101011101" when "0010100", -- t[20] = 861
         "01101000111" when "0010101", -- t[21] = 839
         "01100110001" when "0010110", -- t[22] = 817
         "01100011101" when "0010111", -- t[23] = 797
         "01100001001" when "0011000", -- t[24] = 777
         "01011110110" when "0011001", -- t[25] = 758
         "01011100100" when "0011010", -- t[26] = 740
         "01011010010" when "0011011", -- t[27] = 722
         "01011000001" when "0011100", -- t[28] = 705
         "01010110000" when "0011101", -- t[29] = 688
         "01010100000" when "0011110", -- t[30] = 672
         "01010010001" when "0011111", -- t[31] = 657
         "01010000010" when "0100000", -- t[32] = 642
         "01001110011" when "0100001", -- t[33] = 627
         "01001100101" when "0100010", -- t[34] = 613
         "01001010111" when "0100011", -- t[35] = 599
         "01001001010" when "0100100", -- t[36] = 586
         "01000111110" when "0100101", -- t[37] = 574
         "01000110001" when "0100110", -- t[38] = 561
         "01000100101" when "0100111", -- t[39] = 549
         "01000011010" when "0101000", -- t[40] = 538
         "01000001110" when "0101001", -- t[41] = 526
         "01000000011" when "0101010", -- t[42] = 515
         "00111111001" when "0101011", -- t[43] = 505
         "00111101110" when "0101100", -- t[44] = 494
         "00111100100" when "0101101", -- t[45] = 484
         "00111011011" when "0101110", -- t[46] = 475
         "00111010001" when "0101111", -- t[47] = 465
         "00111001000" when "0110000", -- t[48] = 456
         "00110111111" when "0110001", -- t[49] = 447
         "00110110110" when "0110010", -- t[50] = 438
         "00110101110" when "0110011", -- t[51] = 430
         "00110100110" when "0110100", -- t[52] = 422
         "00110011110" when "0110101", -- t[53] = 414
         "00110010110" when "0110110", -- t[54] = 406
         "00110001110" when "0110111", -- t[55] = 398
         "00110000111" when "0111000", -- t[56] = 391
         "00110000000" when "0111001", -- t[57] = 384
         "00101111001" when "0111010", -- t[58] = 377
         "00101110010" when "0111011", -- t[59] = 370
         "00101101011" when "0111100", -- t[60] = 363
         "00101100101" when "0111101", -- t[61] = 357
         "00101011111" when "0111110", -- t[62] = 351
         "00101011000" when "0111111", -- t[63] = 344
         "00101010010" when "1000000", -- t[64] = 338
         "00101001101" when "1000001", -- t[65] = 333
         "00101000111" when "1000010", -- t[66] = 327
         "00101000001" when "1000011", -- t[67] = 321
         "00100111100" when "1000100", -- t[68] = 316
         "00100110110" when "1000101", -- t[69] = 310
         "00100110001" when "1000110", -- t[70] = 305
         "00100101100" when "1000111", -- t[71] = 300
         "00100100111" when "1001000", -- t[72] = 295
         "00100100010" when "1001001", -- t[73] = 290
         "00100011110" when "1001010", -- t[74] = 286
         "00100011001" when "1001011", -- t[75] = 281
         "00100010101" when "1001100", -- t[76] = 277
         "00100010000" when "1001101", -- t[77] = 272
         "00100001100" when "1001110", -- t[78] = 268
         "00100001000" when "1001111", -- t[79] = 264
         "00100000100" when "1010000", -- t[80] = 260
         "00100000000" when "1010001", -- t[81] = 256
         "00011111100" when "1010010", -- t[82] = 252
         "00011111000" when "1010011", -- t[83] = 248
         "00011110100" when "1010100", -- t[84] = 244
         "00011110000" when "1010101", -- t[85] = 240
         "00011101101" when "1010110", -- t[86] = 237
         "00011101001" when "1010111", -- t[87] = 233
         "00011100110" when "1011000", -- t[88] = 230
         "00011100010" when "1011001", -- t[89] = 226
         "00011011111" when "1011010", -- t[90] = 223
         "00011011100" when "1011011", -- t[91] = 220
         "00011011001" when "1011100", -- t[92] = 217
         "00011010110" when "1011101", -- t[93] = 214
         "00011010010" when "1011110", -- t[94] = 210
         "00011001111" when "1011111", -- t[95] = 207
         "00011001101" when "1100000", -- t[96] = 205
         "00011001010" when "1100001", -- t[97] = 202
         "00011000111" when "1100010", -- t[98] = 199
         "00011000100" when "1100011", -- t[99] = 196
         "00011000001" when "1100100", -- t[100] = 193
         "00010111111" when "1100101", -- t[101] = 191
         "00010111100" when "1100110", -- t[102] = 188
         "00010111010" when "1100111", -- t[103] = 186
         "00010110111" when "1101000", -- t[104] = 183
         "00010110101" when "1101001", -- t[105] = 181
         "00010110010" when "1101010", -- t[106] = 178
         "00010110000" when "1101011", -- t[107] = 176
         "00010101110" when "1101100", -- t[108] = 174
         "00010101011" when "1101101", -- t[109] = 171
         "00010101001" when "1101110", -- t[110] = 169
         "00010100111" when "1101111", -- t[111] = 167
         "00010100101" when "1110000", -- t[112] = 165
         "00010100011" when "1110001", -- t[113] = 163
         "00010100000" when "1110010", -- t[114] = 160
         "00010011110" when "1110011", -- t[115] = 158
         "00010011100" when "1110100", -- t[116] = 156
         "00010011010" when "1110101", -- t[117] = 154
         "00010011001" when "1110110", -- t[118] = 153
         "00010010111" when "1110111", -- t[119] = 151
         "00010010101" when "1111000", -- t[120] = 149
         "00010010011" when "1111001", -- t[121] = 147
         "00010010001" when "1111010", -- t[122] = 145
         "00010001111" when "1111011", -- t[123] = 143
         "00010001110" when "1111100", -- t[124] = 142
         "00010001100" when "1111101", -- t[125] = 140
         "00010001010" when "1111110", -- t[126] = 138
         "00010001001" when "1111111", -- t[127] = 137
         "-----------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_2.
-- Decomposition:
--   alpha_2,2 = 3; sigma'_2,2 = 3; wO_2,2 = 2.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t2_t2 is
  port ( a : in  std_logic_vector(2 downto 0);
         s : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of fp_log_log_23_t2_t2 is
  signal x : std_logic_vector(5 downto 0);
begin
  x <= a & s;

  with x select
    r <= "00" when "000000", -- t[0] = 0
         "00" when "000001", -- t[1] = 0
         "00" when "000010", -- t[2] = 0
         "01" when "000011", -- t[3] = 1
         "01" when "000100", -- t[4] = 1
         "01" when "000101", -- t[5] = 1
         "10" when "000110", -- t[6] = 2
         "10" when "000111", -- t[7] = 2
         "00" when "001000", -- t[8] = 0
         "00" when "001001", -- t[9] = 0
         "00" when "001010", -- t[10] = 0
         "00" when "001011", -- t[11] = 0
         "00" when "001100", -- t[12] = 0
         "01" when "001101", -- t[13] = 1
         "01" when "001110", -- t[14] = 1
         "01" when "001111", -- t[15] = 1
         "00" when "010000", -- t[16] = 0
         "00" when "010001", -- t[17] = 0
         "00" when "010010", -- t[18] = 0
         "00" when "010011", -- t[19] = 0
         "00" when "010100", -- t[20] = 0
         "00" when "010101", -- t[21] = 0
         "00" when "010110", -- t[22] = 0
         "01" when "010111", -- t[23] = 1
         "00" when "011000", -- t[24] = 0
         "00" when "011001", -- t[25] = 0
         "00" when "011010", -- t[26] = 0
         "00" when "011011", -- t[27] = 0
         "00" when "011100", -- t[28] = 0
         "00" when "011101", -- t[29] = 0
         "00" when "011110", -- t[30] = 0
         "00" when "011111", -- t[31] = 0
         "00" when "100000", -- t[32] = 0
         "00" when "100001", -- t[33] = 0
         "00" when "100010", -- t[34] = 0
         "00" when "100011", -- t[35] = 0
         "00" when "100100", -- t[36] = 0
         "00" when "100101", -- t[37] = 0
         "00" when "100110", -- t[38] = 0
         "00" when "100111", -- t[39] = 0
         "00" when "101000", -- t[40] = 0
         "00" when "101001", -- t[41] = 0
         "00" when "101010", -- t[42] = 0
         "00" when "101011", -- t[43] = 0
         "00" when "101100", -- t[44] = 0
         "00" when "101101", -- t[45] = 0
         "00" when "101110", -- t[46] = 0
         "00" when "101111", -- t[47] = 0
         "00" when "110000", -- t[48] = 0
         "00" when "110001", -- t[49] = 0
         "00" when "110010", -- t[50] = 0
         "00" when "110011", -- t[51] = 0
         "00" when "110100", -- t[52] = 0
         "00" when "110101", -- t[53] = 0
         "00" when "110110", -- t[54] = 0
         "00" when "110111", -- t[55] = 0
         "00" when "111000", -- t[56] = 0
         "00" when "111001", -- t[57] = 0
         "00" when "111010", -- t[58] = 0
         "00" when "111011", -- t[59] = 0
         "00" when "111100", -- t[60] = 0
         "00" when "111101", -- t[61] = 0
         "00" when "111110", -- t[62] = 0
         "00" when "111111", -- t[63] = 0
         "--" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 7; beta_2 = 10; lambda_2 = 12;  m_2 = 2;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 7; rho_2,1 = 0; sigma_2,1 = 8; wO_2,1 = 11;
--   Q_2,2 (ROM):  alpha_2,2 = 3; rho_2,2 = 8; sigma_2,2 = 4; wO_2,2 = 2.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23_t2 is
  port ( a : in  std_logic_vector(6 downto 0);
         b : in  std_logic_vector(9 downto 0);
         r : out std_logic_vector(27 downto 0) );
end entity;

architecture arch of fp_log_log_23_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(8 downto 0);
  signal s      : std_logic_vector(11 downto 0);
  component fp_log_log_23_t2_pow is
    port ( x : in  std_logic_vector(8 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  signal a_1    : std_logic_vector(6 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(6 downto 0);
  signal k_1    : std_logic_vector(10 downto 0);
  signal r0_1   : std_logic_vector(19 downto 0);
  signal r_1    : std_logic_vector(27 downto 0);
  component fp_log_log_23_t2_t1 is
    port ( a : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  signal a_2    : std_logic_vector(2 downto 0);
  signal sign_2 : std_logic;
  signal s_2    : std_logic_vector(2 downto 0);
  signal r0_2   : std_logic_vector(1 downto 0);
  signal r_2    : std_logic_vector(27 downto 0);
  component fp_log_log_23_t2_t2 is
    port ( a : in  std_logic_vector(2 downto 0);
           s : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;
begin
  sign <= not b(9);
  b0 <= b(8 downto 0) xor (8 downto 0 => sign);

  pow : fp_log_log_23_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(6 downto 0);
  sign_1 <= not s(11);
  s_1 <= s(10 downto 4) xor (10 downto 4 => sign_1);
  t_1 : fp_log_log_23_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(10 downto 0) <=
    r0_1(19 downto 9) xor (19 downto 9 => ((sign_1)));
  r_1(27 downto 11) <= (27 downto 11 => ((sign_1)));

  a_2 <= a(6 downto 4);
  sign_2 <= not s(3);
  s_2 <= s(2 downto 0) xor (2 downto 0 => sign_2);
  t_2 : fp_log_log_23_t2_t2
    port map ( a => a_2,
               s => s_2,
               r => r0_2 );
  r_2(1 downto 0) <=
    r0_2 xor (1 downto 0 => ((sign_2)));
  r_2(27 downto 2) <= (27 downto 2 => ((sign_2)));

  r <= r_1 + r_2;
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_23 is
  port ( x : in  std_logic_vector(22 downto 0);
         r : out std_logic_vector(27 downto 0) );
end entity;

architecture arch of fp_log_log_23 is
  signal a_0 : std_logic_vector(7 downto 0);
  signal r_0 : std_logic_vector(27 downto 0);
  component fp_log_log_23_t0 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(27 downto 0) );
  end component;

  signal a_1 : std_logic_vector(7 downto 0);
  signal b_1 : std_logic_vector(14 downto 0);
  signal r_1 : std_logic_vector(27 downto 0);
  component fp_log_log_23_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           b : in  std_logic_vector(14 downto 0);
           r : out std_logic_vector(27 downto 0) );
  end component;

  signal a_2 : std_logic_vector(6 downto 0);
  signal b_2 : std_logic_vector(9 downto 0);
  signal r_2 : std_logic_vector(27 downto 0);
  component fp_log_log_23_t2 is
    port ( a : in  std_logic_vector(6 downto 0);
           b : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(27 downto 0) );
  end component;

begin
  a_0 <= x(22 downto 15);
  t_0 : fp_log_log_23_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(22 downto 15);
  b_1 <= x(14 downto 0);
  t_1 : fp_log_log_23_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(22 downto 16);
  b_2 <= x(14 downto 5);
  t_2 : fp_log_log_23_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  r <= r_0 + r_1 + r_2;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- HOTBM instance for function log(x+1/2)/(x-1/2).
-- wI = 24; wO = 24.
-- Order-3 polynomial approximation.
-- Decomposition:
--   alpha = 8; beta = 16;
--   T_0 (ROM):     alpha_0 = 8; beta_0 = 0;
--   T_1 (PowMult): alpha_1 = 8; beta_1 = 16;
--   T_2 (PowMult): alpha_2 = 8; beta_2 = 12;
--   T_3 (ROM):     alpha_3 = 2; beta_3 = 3.
-- Guard bits: g = 4.
-- Command line: logfp 24 24 3   rom 8 0   pm 8 16  ah 16 16 16  1 0  8 16 0   pm 8 12  ah 12 18 9  1 0  8 9 0   rom 2 3


--------------------------------------------------------------------------------
-- TermROM instance for order-0 term.
-- Decomposition:
--   alpha_0 = 8; beta_0 = 0; wO_0 = 29.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t0 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(28 downto 0) );
end entity;

architecture arch of fp_log_log_24_t0 is
  signal x0   : std_logic_vector(7 downto 0);
  signal r0   : std_logic_vector(28 downto 0);
begin
  x0 <= a;

  with x0 select
    r0 <= "10110001001000111011101110111" when "00000000", -- t[0] = 371488631
          "10110000100010000010011111011" when "00000001", -- t[1] = 370214139
          "10101111111011100001010110101" when "00000010", -- t[2] = 368951989
          "10101111010101010111111010111" when "00000011", -- t[3] = 367701975
          "10101110101111100101110011001" when "00000100", -- t[4] = 366463897
          "10101110001010001010100111000" when "00000101", -- t[5] = 365237560
          "10101101100101000101111110100" when "00000110", -- t[6] = 364022772
          "10101101000000010111100010010" when "00000111", -- t[7] = 362819346
          "10101100011011111110111011110" when "00001000", -- t[8] = 361627102
          "10101011110111111011110100100" when "00001001", -- t[9] = 360445860
          "10101011010100001101110110111" when "00001010", -- t[10] = 359275447
          "10101010110000110100101101100" when "00001011", -- t[11] = 358115692
          "10101010001101110000000011101" when "00001100", -- t[12] = 356966429
          "10101001101010111111100101001" when "00001101", -- t[13] = 355827497
          "10101001001000100010111101110" when "00001110", -- t[14] = 354698734
          "10101000100110011001111010100" when "00001111", -- t[15] = 353579988
          "10101000000100100100001000000" when "00010000", -- t[16] = 352471104
          "10100111100011000001010011110" when "00010001", -- t[17] = 351371934
          "10100111000001110001001011110" when "00010010", -- t[18] = 350282334
          "10100110100000110011011101111" when "00010011", -- t[19] = 349202159
          "10100110000000000111111001000" when "00010100", -- t[20] = 348131272
          "10100101011111101110001011111" when "00010101", -- t[21] = 347069535
          "10100100111111100110000101110" when "00010110", -- t[22] = 346016814
          "10100100011111101111010110011" when "00010111", -- t[23] = 344972979
          "10100100000000001001101101110" when "00011000", -- t[24] = 343937902
          "10100011100000110100111100001" when "00011001", -- t[25] = 342911457
          "10100011000001110000110010001" when "00011010", -- t[26] = 341893521
          "10100010100010111101000000110" when "00011011", -- t[27] = 340883974
          "10100010000100011001011001001" when "00011100", -- t[28] = 339882697
          "10100001100110000101101101000" when "00011101", -- t[29] = 338889576
          "10100001001000000001101110000" when "00011110", -- t[30] = 337904496
          "10100000101010001101001110011" when "00011111", -- t[31] = 336927347
          "10100000001100101000000000011" when "00100000", -- t[32] = 335958019
          "10011111101111010001110110110" when "00100001", -- t[33] = 334996406
          "10011111010010001010100100011" when "00100010", -- t[34] = 334042403
          "10011110110101010001111100100" when "00100011", -- t[35] = 333095908
          "10011110011000100111110010011" when "00100100", -- t[36] = 332156819
          "10011101111100001011111001111" when "00100101", -- t[37] = 331225039
          "10011101011111111110000110101" when "00100110", -- t[38] = 330300469
          "10011101000011111110001100111" when "00100111", -- t[39] = 329383015
          "10011100101000001100000001001" when "00101000", -- t[40] = 328472585
          "10011100001100100111010111101" when "00101001", -- t[41] = 327569085
          "10011011110001010000000101010" when "00101010", -- t[42] = 326672426
          "10011011010110000101111111001" when "00101011", -- t[43] = 325782521
          "10011010111011001000111010010" when "00101100", -- t[44] = 324899282
          "10011010100000011000101100000" when "00101101", -- t[45] = 324022624
          "10011010000101110101001010001" when "00101110", -- t[46] = 323152465
          "10011001101011011110001010001" when "00101111", -- t[47] = 322288721
          "10011001010001010011100010001" when "00110000", -- t[48] = 321431313
          "10011000110111010101001000010" when "00110001", -- t[49] = 320580162
          "10011000011101100010110010110" when "00110010", -- t[50] = 319735190
          "10011000000011111100011000001" when "00110011", -- t[51] = 318896321
          "10010111101010100001101110111" when "00110100", -- t[52] = 318063479
          "10010111010001010010101110000" when "00110101", -- t[53] = 317236592
          "10010110111000001111001100010" when "00110110", -- t[54] = 316415586
          "10010110011111010111000000111" when "00110111", -- t[55] = 315600391
          "10010110000110101010000011001" when "00111000", -- t[56] = 314790937
          "10010101101110001000001010100" when "00111001", -- t[57] = 313987156
          "10010101010101110001001110011" when "00111010", -- t[58] = 313188979
          "10010100111101100101000110100" when "00111011", -- t[59] = 312396340
          "10010100100101100011101010111" when "00111100", -- t[60] = 311609175
          "10010100001101101100110011010" when "00111101", -- t[61] = 310827418
          "10010011110110000000011000000" when "00111110", -- t[62] = 310051008
          "10010011011110011110010001001" when "00111111", -- t[63] = 309279881
          "10010011000111000110010111010" when "01000000", -- t[64] = 308513978
          "10010010101111111000100010101" when "01000001", -- t[65] = 307753237
          "10010010011000110100101100000" when "01000010", -- t[66] = 306997600
          "10010010000001111010101100001" when "01000011", -- t[67] = 306247009
          "10010001101011001010011011111" when "01000100", -- t[68] = 305501407
          "10010001010100100011110100001" when "01000101", -- t[69] = 304760737
          "10010000111110000110101110001" when "01000110", -- t[70] = 304024945
          "10010000100111110011000010111" when "01000111", -- t[71] = 303293975
          "10010000010001101000101011110" when "01001000", -- t[72] = 302567774
          "10001111111011100111100010010" when "01001001", -- t[73] = 301846290
          "10001111100101101111011111111" when "01001010", -- t[74] = 301129471
          "10001111010000000000011110001" when "01001011", -- t[75] = 300417265
          "10001110111010011010010110110" when "01001100", -- t[76] = 299709622
          "10001110100100111101000011101" when "01001101", -- t[77] = 299006493
          "10001110001111101000011110101" when "01001110", -- t[78] = 298307829
          "10001101111010011100100001110" when "01001111", -- t[79] = 297613582
          "10001101100101011001000111001" when "01010000", -- t[80] = 296923705
          "10001101010000011110001000111" when "01010001", -- t[81] = 296238151
          "10001100111011101011100001011" when "01010010", -- t[82] = 295556875
          "10001100100111000001001010111" when "01010011", -- t[83] = 294879831
          "10001100010010011110111111110" when "01010100", -- t[84] = 294206974
          "10001011111110000100111010110" when "01010101", -- t[85] = 293538262
          "10001011101001110010110110010" when "01010110", -- t[86] = 292873650
          "10001011010101101000101101001" when "01010111", -- t[87] = 292213097
          "10001011000001100110011010000" when "01011000", -- t[88] = 291556560
          "10001010101101101011110111111" when "01011001", -- t[89] = 290903999
          "10001010011001111001000001011" when "01011010", -- t[90] = 290255371
          "10001010000110001101110001111" when "01011011", -- t[91] = 289610639
          "10001001110010101010000100001" when "01011100", -- t[92] = 288969761
          "10001001011111001101110011011" when "01011101", -- t[93] = 288332699
          "10001001001011111000111010111" when "01011110", -- t[94] = 287699415
          "10001000111000101011010101110" when "01011111", -- t[95] = 287069870
          "10001000100101100100111111100" when "01100000", -- t[96] = 286444028
          "10001000010010100101110011100" when "01100001", -- t[97] = 285821852
          "10000111111111101101101101001" when "01100010", -- t[98] = 285203305
          "10000111101100111100101000000" when "01100011", -- t[99] = 284588352
          "10000111011010010010011111101" when "01100100", -- t[100] = 283976957
          "10000111000111101111001111110" when "01100101", -- t[101] = 283369086
          "10000110110101010010110100001" when "01100110", -- t[102] = 282764705
          "10000110100010111101001000011" when "01100111", -- t[103] = 282163779
          "10000110010000101110001000100" when "01101000", -- t[104] = 281566276
          "10000101111110100101110000010" when "01101001", -- t[105] = 280972162
          "10000101101100100011111011101" when "01101010", -- t[106] = 280381405
          "10000101011010101000100110110" when "01101011", -- t[107] = 279793974
          "10000101001000110011101101100" when "01101100", -- t[108] = 279209836
          "10000100110111000101001100000" when "01101101", -- t[109] = 278628960
          "10000100100101011100111110100" when "01101110", -- t[110] = 278051316
          "10000100010011111011000001010" when "01101111", -- t[111] = 277476874
          "10000100000010011111010000011" when "01110000", -- t[112] = 276905603
          "10000011110001001001101000010" when "01110001", -- t[113] = 276337474
          "10000011011111111010000101010" when "01110010", -- t[114] = 275772458
          "10000011001110110000100011110" when "01110011", -- t[115] = 275210526
          "10000010111101101101000000010" when "01110100", -- t[116] = 274651650
          "10000010101100101111010111010" when "01110101", -- t[117] = 274095802
          "10000010011011110111100101010" when "01110110", -- t[118] = 273542954
          "10000010001011000101100110111" when "01110111", -- t[119] = 272993079
          "10000001111010011001011000110" when "01111000", -- t[120] = 272446150
          "10000001101001110010110111100" when "01111001", -- t[121] = 271902140
          "10000001011001010010000000000" when "01111010", -- t[122] = 271361024
          "10000001001000110110101110111" when "01111011", -- t[123] = 270822775
          "10000000111000100001000001000" when "01111100", -- t[124] = 270287368
          "10000000101000010000110011010" when "01111101", -- t[125] = 269754778
          "10000000011000000110000010011" when "01111110", -- t[126] = 269224979
          "10000000001000000000101011011" when "01111111", -- t[127] = 268697947
          "01111111111000000000101011010" when "10000000", -- t[128] = 268173658
          "01111111101000000101111111000" when "10000001", -- t[129] = 267652088
          "01111111011000010000100011101" when "10000010", -- t[130] = 267133213
          "01111111001000100000010110001" when "10000011", -- t[131] = 266617009
          "01111110111000110101010011110" when "10000100", -- t[132] = 266103454
          "01111110101001001111011001100" when "10000101", -- t[133] = 265592524
          "01111110011001101110100100110" when "10000110", -- t[134] = 265084198
          "01111110001010010010110010100" when "10000111", -- t[135] = 264578452
          "01111101111010111100000000010" when "10001000", -- t[136] = 264075266
          "01111101101011101010001011000" when "10001001", -- t[137] = 263574616
          "01111101011100011101010000010" when "10001010", -- t[138] = 263076482
          "01111101001101010101001101010" when "10001011", -- t[139] = 262580842
          "01111100111110010001111111011" when "10001100", -- t[140] = 262087675
          "01111100101111010011100100001" when "10001101", -- t[141] = 261596961
          "01111100100000011001111001000" when "10001110", -- t[142] = 261108680
          "01111100010001100100111011010" when "10001111", -- t[143] = 260622810
          "01111100000010110100101000100" when "10010000", -- t[144] = 260139332
          "01111011110100001000111110010" when "10010001", -- t[145] = 259658226
          "01111011100101100001111010001" when "10010010", -- t[146] = 259179473
          "01111011010110111111011001101" when "10010011", -- t[147] = 258703053
          "01111011001000100001011010100" when "10010100", -- t[148] = 258228948
          "01111010111010000111111010001" when "10010101", -- t[149] = 257757137
          "01111010101011110010110110100" when "10010110", -- t[150] = 257287604
          "01111010011101100010001101001" when "10010111", -- t[151] = 256820329
          "01111010001111010101111011110" when "10011000", -- t[152] = 256355294
          "01111010000001001110000000001" when "10011001", -- t[153] = 255892481
          "01111001110011001010011000000" when "10011010", -- t[154] = 255431872
          "01111001100101001011000001010" when "10011011", -- t[155] = 254973450
          "01111001010111001111111001101" when "10011100", -- t[156] = 254517197
          "01111001001001011000111111000" when "10011101", -- t[157] = 254063096
          "01111000111011100110001111010" when "10011110", -- t[158] = 253611130
          "01111000101101110111101000011" when "10011111", -- t[159] = 253161283
          "01111000100000001101001000001" when "10100000", -- t[160] = 252713537
          "01111000010010100110101100100" when "10100001", -- t[161] = 252267876
          "01111000000101000100010011100" when "10100010", -- t[162] = 251824284
          "01110111110111100101111011001" when "10100011", -- t[163] = 251382745
          "01110111101010001011100001010" when "10100100", -- t[164] = 250943242
          "01110111011100110101000100001" when "10100101", -- t[165] = 250505761
          "01110111001111100010100001101" when "10100110", -- t[166] = 250070285
          "01110111000010010011111000000" when "10100111", -- t[167] = 249636800
          "01110110110101001001000101001" when "10101000", -- t[168] = 249205289
          "01110110101000000010000111010" when "10101001", -- t[169] = 248775738
          "01110110011010111110111100101" when "10101010", -- t[170] = 248348133
          "01110110001101111111100011001" when "10101011", -- t[171] = 247922457
          "01110110000001000011111001001" when "10101100", -- t[172] = 247498697
          "01110101110100001011111100110" when "10101101", -- t[173] = 247076838
          "01110101100111010111101100010" when "10101110", -- t[174] = 246656866
          "01110101011010100111000101111" when "10101111", -- t[175] = 246238767
          "01110101001101111010000111111" when "10110000", -- t[176] = 245822527
          "01110101000001010000110000100" when "10110001", -- t[177] = 245408132
          "01110100110100101010111110000" when "10110010", -- t[178] = 244995568
          "01110100101000001000101110110" when "10110011", -- t[179] = 244584822
          "01110100011011101010000001000" when "10110100", -- t[180] = 244175880
          "01110100001111001110110011010" when "10110101", -- t[181] = 243768730
          "01110100000010110111000011101" when "10110110", -- t[182] = 243363357
          "01110011110110100010110000110" when "10110111", -- t[183] = 242959750
          "01110011101010010001111000111" when "10111000", -- t[184] = 242557895
          "01110011011110000100011010011" when "10111001", -- t[185] = 242157779
          "01110011010001111010010011110" when "10111010", -- t[186] = 241759390
          "01110011000101110011100011011" when "10111011", -- t[187] = 241362715
          "01110010111001110000000111111" when "10111100", -- t[188] = 240967743
          "01110010101101101111111111100" when "10111101", -- t[189] = 240574460
          "01110010100001110011001001000" when "10111110", -- t[190] = 240182856
          "01110010010101111001100010101" when "10111111", -- t[191] = 239792917
          "01110010001010000011001011000" when "11000000", -- t[192] = 239404632
          "01110001111110010000000000101" when "11000001", -- t[193] = 239017989
          "01110001110010100000000010001" when "11000010", -- t[194] = 238632977
          "01110001100110110011001110001" when "11000011", -- t[195] = 238249585
          "01110001011011001001100011000" when "11000100", -- t[196] = 237867800
          "01110001001111100010111111100" when "11000101", -- t[197] = 237487612
          "01110001000011111111100010001" when "11000110", -- t[198] = 237109009
          "01110000111000011111001001100" when "11000111", -- t[199] = 236731980
          "01110000101101000001110100011" when "11001000", -- t[200] = 236356515
          "01110000100001100111100001011" when "11001001", -- t[201] = 235982603
          "01110000010110010000001111000" when "11001010", -- t[202] = 235610232
          "01110000001010111011111100001" when "11001011", -- t[203] = 235239393
          "01101111111111101010100111011" when "11001100", -- t[204] = 234870075
          "01101111110100011100001111011" when "11001101", -- t[205] = 234502267
          "01101111101001010000110010111" when "11001110", -- t[206] = 234135959
          "01101111011110001000010000101" when "11001111", -- t[207] = 233771141
          "01101111010011000010100111010" when "11010000", -- t[208] = 233407802
          "01101111000111111111110101110" when "11010001", -- t[209] = 233045934
          "01101110111100111111111010101" when "11010010", -- t[210] = 232685525
          "01101110110010000010110100110" when "11010011", -- t[211] = 232326566
          "01101110100111001000100011000" when "11010100", -- t[212] = 231969048
          "01101110011100010001000100000" when "11010101", -- t[213] = 231612960
          "01101110010001011100010110101" when "11010110", -- t[214] = 231258293
          "01101110000110101010011001110" when "11010111", -- t[215] = 230905038
          "01101101111011111011001100001" when "11011000", -- t[216] = 230553185
          "01101101110001001110101100110" when "11011001", -- t[217] = 230202726
          "01101101100110100100111010010" when "11011010", -- t[218] = 229853650
          "01101101011011111101110011100" when "11011011", -- t[219] = 229505948
          "01101101010001011001010111101" when "11011100", -- t[220] = 229159613
          "01101101000110110111100101010" when "11011101", -- t[221] = 228814634
          "01101100111100011000011011011" when "11011110", -- t[222] = 228471003
          "01101100110001111011111000111" when "11011111", -- t[223] = 228128711
          "01101100100111100001111100101" when "11100000", -- t[224] = 227787749
          "01101100011101001010100101101" when "11100001", -- t[225] = 227448109
          "01101100010010110101110010111" when "11100010", -- t[226] = 227109783
          "01101100001000100011100011001" when "11100011", -- t[227] = 226772761
          "01101011111110010011110101100" when "11100100", -- t[228] = 226437036
          "01101011110100000110101000111" when "11100101", -- t[229] = 226102599
          "01101011101001111011111100001" when "11100110", -- t[230] = 225769441
          "01101011011111110011101110100" when "11100111", -- t[231] = 225437556
          "01101011010101101101111110110" when "11101000", -- t[232] = 225106934
          "01101011001011101010101011111" when "11101001", -- t[233] = 224777567
          "01101011000001101001110101001" when "11101010", -- t[234] = 224449449
          "01101010110111101011011001010" when "11101011", -- t[235] = 224122570
          "01101010101101101111010111011" when "11101100", -- t[236] = 223796923
          "01101010100011110101101110101" when "11101101", -- t[237] = 223472501
          "01101010011001111110011101111" when "11101110", -- t[238] = 223149295
          "01101010010000001001100100010" when "11101111", -- t[239] = 222827298
          "01101010000110010111000000111" when "11110000", -- t[240] = 222506503
          "01101001111100100110110010101" when "11110001", -- t[241] = 222186901
          "01101001110010111000111000111" when "11110010", -- t[242] = 221868487
          "01101001101001001101010010100" when "11110011", -- t[243] = 221551252
          "01101001011111100011111110100" when "11110100", -- t[244] = 221235188
          "01101001010101111100111100010" when "11110101", -- t[245] = 220920290
          "01101001001100011000001010110" when "11110110", -- t[246] = 220606550
          "01101001000010110101101001000" when "11110111", -- t[247] = 220293960
          "01101000111001010101010110001" when "11111000", -- t[248] = 219982513
          "01101000101111110111010001100" when "11111001", -- t[249] = 219672204
          "01101000100110011011011010000" when "11111010", -- t[250] = 219363024
          "01101000011101000001101110111" when "11111011", -- t[251] = 219054967
          "01101000010011101010001111010" when "11111100", -- t[252] = 218748026
          "01101000001010010100111010011" when "11111101", -- t[253] = 218442195
          "01101000000001000001101111010" when "11111110", -- t[254] = 218137466
          "01100111110111110000101101001" when "11111111", -- t[255] = 217833833
          "-----------------------------" when others;

  r(28 downto 0) <= r0;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-1 powering unit.
-- Decomposition:
--   beta_1 = 16; mu_1 = 16; lambda_1 = 16.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t1_pow is
  port ( x : in  std_logic_vector(14 downto 0);
         r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of fp_log_log_24_t1_pow is
  signal pp0 : std_logic_vector(14 downto 0);
  signal r0 : std_logic_vector(14 downto 0);
begin
  pp0(14) <= x(14);

  pp0(13) <= x(13);

  pp0(12) <= x(12);

  pp0(11) <= x(11);

  pp0(10) <= x(10);

  pp0(9) <= x(9);

  pp0(8) <= x(8);

  pp0(7) <= x(7);

  pp0(6) <= x(6);

  pp0(5) <= x(5);

  pp0(4) <= x(4);

  pp0(3) <= x(3);

  pp0(2) <= x(2);

  pp0(1) <= x(1);

  pp0(0) <= x(0);

  r0 <= pp0;
  r <= "1" & r0(14 downto 0);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-1 term Q_1.
-- Decomposition:
--   alpha_1,1 = 8; wO_1,1 = 21.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t1_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(20 downto 0) );
end entity;

architecture arch of fp_log_log_24_t1_t1 is
  signal x : std_logic_vector(7 downto 0);
begin
  x <= a;

  with x select
    r <= "100111000101011011100" when "00000000", -- t[0] = 1280732
         "100110101101000111110" when "00000001", -- t[1] = 1268286
         "100110010101001110000" when "00000010", -- t[2] = 1256048
         "100101111101101101101" when "00000011", -- t[3] = 1244013
         "100101100110100110000" when "00000100", -- t[4] = 1232176
         "100101001111110110011" when "00000101", -- t[5] = 1220531
         "100100111001011110100" when "00000110", -- t[6] = 1209076
         "100100100011011101101" when "00000111", -- t[7] = 1197805
         "100100001101110011010" when "00001000", -- t[8] = 1186714
         "100011111000011110111" when "00001001", -- t[9] = 1175799
         "100011100011100000000" when "00001010", -- t[10] = 1165056
         "100011001110110110001" when "00001011", -- t[11] = 1154481
         "100010111010100000111" when "00001100", -- t[12] = 1144071
         "100010100110011111101" when "00001101", -- t[13] = 1133821
         "100010010010110010001" when "00001110", -- t[14] = 1123729
         "100001111111010111110" when "00001111", -- t[15] = 1113790
         "100001101100010000010" when "00010000", -- t[16] = 1104002
         "100001011001011011001" when "00010001", -- t[17] = 1094361
         "100001000110111000000" when "00010010", -- t[18] = 1084864
         "100000110100100110100" when "00010011", -- t[19] = 1075508
         "100000100010100110010" when "00010100", -- t[20] = 1066290
         "100000010000110110111" when "00010101", -- t[21] = 1057207
         "011111111111011000000" when "00010110", -- t[22] = 1048256
         "011111101110001001011" when "00010111", -- t[23] = 1039435
         "011111011101001010100" when "00011000", -- t[24] = 1030740
         "011111001100011011010" when "00011001", -- t[25] = 1022170
         "011110111011111011010" when "00011010", -- t[26] = 1013722
         "011110101011101010000" when "00011011", -- t[27] = 1005392
         "011110011011100111100" when "00011100", -- t[28] = 997180
         "011110001011110011010" when "00011101", -- t[29] = 989082
         "011101111100001101000" when "00011110", -- t[30] = 981096
         "011101101100110100101" when "00011111", -- t[31] = 973221
         "011101011101101001101" when "00100000", -- t[32] = 965453
         "011101001110101011111" when "00100001", -- t[33] = 957791
         "011100111111111011000" when "00100010", -- t[34] = 950232
         "011100110001010110111" when "00100011", -- t[35] = 942775
         "011100100010111111010" when "00100100", -- t[36] = 935418
         "011100010100110011111" when "00100101", -- t[37] = 928159
         "011100000110110100100" when "00100110", -- t[38] = 920996
         "011011111001000000111" when "00100111", -- t[39] = 913927
         "011011101011011000110" when "00101000", -- t[40] = 906950
         "011011011101111100000" when "00101001", -- t[41] = 900064
         "011011010000101010011" when "00101010", -- t[42] = 893267
         "011011000011100011110" when "00101011", -- t[43] = 886558
         "011010110110100111110" when "00101100", -- t[44] = 879934
         "011010101001110110011" when "00101101", -- t[45] = 873395
         "011010011101001111010" when "00101110", -- t[46] = 866938
         "011010010000110010010" when "00101111", -- t[47] = 860562
         "011010000100011111010" when "00110000", -- t[48] = 854266
         "011001111000010110001" when "00110001", -- t[49] = 848049
         "011001101100010110100" when "00110010", -- t[50] = 841908
         "011001100000100000011" when "00110011", -- t[51] = 835843
         "011001010100110011100" when "00110100", -- t[52] = 829852
         "011001001001001111111" when "00110101", -- t[53] = 823935
         "011000111101110101000" when "00110110", -- t[54] = 818088
         "011000110010100011001" when "00110111", -- t[55] = 812313
         "011000100111011001110" when "00111000", -- t[56] = 806606
         "011000011100011001000" when "00111001", -- t[57] = 800968
         "011000010001100000101" when "00111010", -- t[58] = 795397
         "011000000110110000011" when "00111011", -- t[59] = 789891
         "010111111100001000010" when "00111100", -- t[60] = 784450
         "010111110001101000001" when "00111101", -- t[61] = 779073
         "010111100111001111110" when "00111110", -- t[62] = 773758
         "010111011100111111001" when "00111111", -- t[63] = 768505
         "010111010010110110000" when "01000000", -- t[64] = 763312
         "010111001000110100011" when "01000001", -- t[65] = 758179
         "010110111110111010000" when "01000010", -- t[66] = 753104
         "010110110101000110111" when "01000011", -- t[67] = 748087
         "010110101011011010111" when "01000100", -- t[68] = 743127
         "010110100001110101110" when "01000101", -- t[69] = 738222
         "010110011000010111100" when "01000110", -- t[70] = 733372
         "010110001111000000000" when "01000111", -- t[71] = 728576
         "010110000101101111010" when "01001000", -- t[72] = 723834
         "010101111100100100111" when "01001001", -- t[73] = 719143
         "010101110011100001000" when "01001010", -- t[74] = 714504
         "010101101010100011100" when "01001011", -- t[75] = 709916
         "010101100001101100010" when "01001100", -- t[76] = 705378
         "010101011000111011000" when "01001101", -- t[77] = 700888
         "010101010000001111111" when "01001110", -- t[78] = 696447
         "010101000111101010110" when "01001111", -- t[79] = 692054
         "010100111111001011100" when "01010000", -- t[80] = 687708
         "010100110110110010000" when "01010001", -- t[81] = 683408
         "010100101110011110001" when "01010010", -- t[82] = 679153
         "010100100110001111111" when "01010011", -- t[83] = 674943
         "010100011110000111001" when "01010100", -- t[84] = 670777
         "010100010110000011111" when "01010101", -- t[85] = 666655
         "010100001110000101111" when "01010110", -- t[86] = 662575
         "010100000110001101010" when "01010111", -- t[87] = 658538
         "010011111110011001110" when "01011000", -- t[88] = 654542
         "010011110110101011100" when "01011001", -- t[89] = 650588
         "010011101111000010001" when "01011010", -- t[90] = 646673
         "010011100111011101111" when "01011011", -- t[91] = 642799
         "010011011111111110011" when "01011100", -- t[92] = 638963
         "010011011000100011111" when "01011101", -- t[93] = 635167
         "010011010001001110000" when "01011110", -- t[94] = 631408
         "010011001001111100111" when "01011111", -- t[95] = 627687
         "010011000010110000011" when "01100000", -- t[96] = 624003
         "010010111011101000100" when "01100001", -- t[97] = 620356
         "010010110100100101000" when "01100010", -- t[98] = 616744
         "010010101101100110000" when "01100011", -- t[99] = 613168
         "010010100110101011011" when "01100100", -- t[100] = 609627
         "010010011111110101000" when "01100101", -- t[101] = 606120
         "010010011001000011000" when "01100110", -- t[102] = 602648
         "010010010010010101001" when "01100111", -- t[103] = 599209
         "010010001011101011011" when "01101000", -- t[104] = 595803
         "010010000101000101110" when "01101001", -- t[105] = 592430
         "010001111110100100001" when "01101010", -- t[106] = 589089
         "010001111000000110100" when "01101011", -- t[107] = 585780
         "010001110001101100110" when "01101100", -- t[108] = 582502
         "010001101011010110111" when "01101101", -- t[109] = 579255
         "010001100101000100110" when "01101110", -- t[110] = 576038
         "010001011110110110100" when "01101111", -- t[111] = 572852
         "010001011000101011111" when "01110000", -- t[112] = 569695
         "010001010010100101000" when "01110001", -- t[113] = 566568
         "010001001100100001101" when "01110010", -- t[114] = 563469
         "010001000110100001111" when "01110011", -- t[115] = 560399
         "010001000000100101101" when "01110100", -- t[116] = 557357
         "010000111010101100111" when "01110101", -- t[117] = 554343
         "010000110100110111101" when "01110110", -- t[118] = 551357
         "010000101111000101101" when "01110111", -- t[119] = 548397
         "010000101001010111001" when "01111000", -- t[120] = 545465
         "010000100011101011110" when "01111001", -- t[121] = 542558
         "010000011110000011110" when "01111010", -- t[122] = 539678
         "010000011000011111000" when "01111011", -- t[123] = 536824
         "010000010010111101011" when "01111100", -- t[124] = 533995
         "010000001101011110110" when "01111101", -- t[125] = 531190
         "010000001000000011011" when "01111110", -- t[126] = 528411
         "010000000010101011000" when "01111111", -- t[127] = 525656
         "001111111101010101110" when "10000000", -- t[128] = 522926
         "001111111000000011011" when "10000001", -- t[129] = 520219
         "001111110010110100000" when "10000010", -- t[130] = 517536
         "001111101101100111100" when "10000011", -- t[131] = 514876
         "001111101000011101111" when "10000100", -- t[132] = 512239
         "001111100011010111000" when "10000101", -- t[133] = 509624
         "001111011110010011000" when "10000110", -- t[134] = 507032
         "001111011001010001111" when "10000111", -- t[135] = 504463
         "001111010100010011011" when "10001000", -- t[136] = 501915
         "001111001111010111100" when "10001001", -- t[137] = 499388
         "001111001010011110100" when "10001010", -- t[138] = 496884
         "001111000101101000000" when "10001011", -- t[139] = 494400
         "001111000000110100001" when "10001100", -- t[140] = 491937
         "001110111100000010110" when "10001101", -- t[141] = 489494
         "001110110111010100000" when "10001110", -- t[142] = 487072
         "001110110010100111111" when "10001111", -- t[143] = 484671
         "001110101101111110001" when "10010000", -- t[144] = 482289
         "001110101001010110110" when "10010001", -- t[145] = 479926
         "001110100100110001111" when "10010010", -- t[146] = 477583
         "001110100000001111100" when "10010011", -- t[147] = 475260
         "001110011011101111011" when "10010100", -- t[148] = 472955
         "001110010111010001101" when "10010101", -- t[149] = 470669
         "001110010010110110001" when "10010110", -- t[150] = 468401
         "001110001110011101000" when "10010111", -- t[151] = 466152
         "001110001010000110001" when "10011000", -- t[152] = 463921
         "001110000101110001100" when "10011001", -- t[153] = 461708
         "001110000001011111001" when "10011010", -- t[154] = 459513
         "001101111101001110111" when "10011011", -- t[155] = 457335
         "001101111001000000110" when "10011100", -- t[156] = 455174
         "001101110100110100110" when "10011101", -- t[157] = 453030
         "001101110000101011000" when "10011110", -- t[158] = 450904
         "001101101100100011010" when "10011111", -- t[159] = 448794
         "001101101000011101101" when "10100000", -- t[160] = 446701
         "001101100100011010000" when "10100001", -- t[161] = 444624
         "001101100000011000011" when "10100010", -- t[162] = 442563
         "001101011100011000110" when "10100011", -- t[163] = 440518
         "001101011000011011001" when "10100100", -- t[164] = 438489
         "001101010100011111100" when "10100101", -- t[165] = 436476
         "001101010000100101110" when "10100110", -- t[166] = 434478
         "001101001100101110000" when "10100111", -- t[167] = 432496
         "001101001000111000000" when "10101000", -- t[168] = 430528
         "001101000101000100000" when "10101001", -- t[169] = 428576
         "001101000001010001110" when "10101010", -- t[170] = 426638
         "001100111101100001011" when "10101011", -- t[171] = 424715
         "001100111001110010111" when "10101100", -- t[172] = 422807
         "001100110110000110001" when "10101101", -- t[173] = 420913
         "001100110010011011001" when "10101110", -- t[174] = 419033
         "001100101110110001111" when "10101111", -- t[175] = 417167
         "001100101011001010011" when "10110000", -- t[176] = 415315
         "001100100111100100101" when "10110001", -- t[177] = 413477
         "001100100100000000101" when "10110010", -- t[178] = 411653
         "001100100000011110010" when "10110011", -- t[179] = 409842
         "001100011100111101100" when "10110100", -- t[180] = 408044
         "001100011001011110011" when "10110101", -- t[181] = 406259
         "001100010110000001000" when "10110110", -- t[182] = 404488
         "001100010010100101001" when "10110111", -- t[183] = 402729
         "001100001111001010111" when "10111000", -- t[184] = 400983
         "001100001011110010010" when "10111001", -- t[185] = 399250
         "001100001000011011010" when "10111010", -- t[186] = 397530
         "001100000101000101101" when "10111011", -- t[187] = 395821
         "001100000001110001101" when "10111100", -- t[188] = 394125
         "001011111110011111010" when "10111101", -- t[189] = 392442
         "001011111011001110010" when "10111110", -- t[190] = 390770
         "001011110111111110110" when "10111111", -- t[191] = 389110
         "001011110100110000110" when "11000000", -- t[192] = 387462
         "001011110001100100001" when "11000001", -- t[193] = 385825
         "001011101110011001000" when "11000010", -- t[194] = 384200
         "001011101011001111011" when "11000011", -- t[195] = 382587
         "001011101000000111001" when "11000100", -- t[196] = 380985
         "001011100101000000010" when "11000101", -- t[197] = 379394
         "001011100001111010110" when "11000110", -- t[198] = 377814
         "001011011110110110101" when "11000111", -- t[199] = 376245
         "001011011011110011111" when "11001000", -- t[200] = 374687
         "001011011000110010100" when "11001001", -- t[201] = 373140
         "001011010101110010011" when "11001010", -- t[202] = 371603
         "001011010010110011101" when "11001011", -- t[203] = 370077
         "001011001111110110001" when "11001100", -- t[204] = 368561
         "001011001100111010000" when "11001101", -- t[205] = 367056
         "001011001001111111001" when "11001110", -- t[206] = 365561
         "001011000111000101101" when "11001111", -- t[207] = 364077
         "001011000100001101010" when "11010000", -- t[208] = 362602
         "001011000001010110001" when "11010001", -- t[209] = 361137
         "001010111110100000010" when "11010010", -- t[210] = 359682
         "001010111011101011101" when "11010011", -- t[211] = 358237
         "001010111000111000010" when "11010100", -- t[212] = 356802
         "001010110110000110000" when "11010101", -- t[213] = 355376
         "001010110011010100111" when "11010110", -- t[214] = 353959
         "001010110000100101000" when "11010111", -- t[215] = 352552
         "001010101101110110011" when "11011000", -- t[216] = 351155
         "001010101011001000110" when "11011001", -- t[217] = 349766
         "001010101000011100011" when "11011010", -- t[218] = 348387
         "001010100101110001001" when "11011011", -- t[219] = 347017
         "001010100011000111000" when "11011100", -- t[220] = 345656
         "001010100000011110000" when "11011101", -- t[221] = 344304
         "001010011101110110000" when "11011110", -- t[222] = 342960
         "001010011011001111001" when "11011111", -- t[223] = 341625
         "001010011000101001011" when "11100000", -- t[224] = 340299
         "001010010110000100110" when "11100001", -- t[225] = 338982
         "001010010011100001001" when "11100010", -- t[226] = 337673
         "001010010000111110100" when "11100011", -- t[227] = 336372
         "001010001110011101000" when "11100100", -- t[228] = 335080
         "001010001011111100100" when "11100101", -- t[229] = 333796
         "001010001001011101000" when "11100110", -- t[230] = 332520
         "001010000110111110100" when "11100111", -- t[231] = 331252
         "001010000100100001001" when "11101000", -- t[232] = 329993
         "001010000010000100101" when "11101001", -- t[233] = 328741
         "001001111111101001001" when "11101010", -- t[234] = 327497
         "001001111101001110110" when "11101011", -- t[235] = 326262
         "001001111010110101001" when "11101100", -- t[236] = 325033
         "001001111000011100101" when "11101101", -- t[237] = 323813
         "001001110110000101000" when "11101110", -- t[238] = 322600
         "001001110011101110011" when "11101111", -- t[239] = 321395
         "001001110001011000101" when "11110000", -- t[240] = 320197
         "001001101111000011111" when "11110001", -- t[241] = 319007
         "001001101100110000000" when "11110010", -- t[242] = 317824
         "001001101010011101000" when "11110011", -- t[243] = 316648
         "001001101000001011000" when "11110100", -- t[244] = 315480
         "001001100101111001110" when "11110101", -- t[245] = 314318
         "001001100011101001100" when "11110110", -- t[246] = 313164
         "001001100001011010001" when "11110111", -- t[247] = 312017
         "001001011111001011101" when "11111000", -- t[248] = 310877
         "001001011100111110000" when "11111001", -- t[249] = 309744
         "001001011010110001001" when "11111010", -- t[250] = 308617
         "001001011000100101010" when "11111011", -- t[251] = 307498
         "001001010110011010001" when "11111100", -- t[252] = 306385
         "001001010100001111111" when "11111101", -- t[253] = 305279
         "001001010010000110011" when "11111110", -- t[254] = 304179
         "001001001111111101111" when "11111111", -- t[255] = 303087
         "---------------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-1 term.
-- Decomposition:
--   alpha_1 = 8; beta_1 = 16; lambda_1 = 16;  m_1 = 1;
--   Pow   (AdHoc);
--   Q_1,1 (Mult): alpha_1,1 = 8; rho_1,1 = 0; sigma_1,1 = 16; wO_1,1 = 21.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         b : in  std_logic_vector(15 downto 0);
         r : out std_logic_vector(28 downto 0) );
end entity;

architecture arch of fp_log_log_24_t1 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(14 downto 0);
  signal s      : std_logic_vector(15 downto 0);
  component fp_log_log_24_t1_pow is
    port ( x : in  std_logic_vector(14 downto 0);
           r : out std_logic_vector(15 downto 0) );
  end component;

  signal a_1    : std_logic_vector(7 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(14 downto 0);
  signal k_1    : std_logic_vector(20 downto 0);
  signal r0_1   : std_logic_vector(37 downto 0);
  signal r_1    : std_logic_vector(28 downto 0);
  component fp_log_log_24_t1_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(20 downto 0) );
  end component;
begin
  sign <= not b(15);
  b0 <= b(14 downto 0) xor (14 downto 0 => sign);

  pow : fp_log_log_24_t1_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(7 downto 0);
  sign_1 <= not s(15);
  s_1 <= s(14 downto 0) xor (14 downto 0 => sign_1);
  t_1 : fp_log_log_24_t1_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(20 downto 0) <=
    r0_1(37 downto 17) xor (37 downto 17 => (not (sign xor sign_1)));
  r_1(28 downto 21) <= (28 downto 21 => (not (sign xor sign_1)));

  r <= r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_fp_log.all;

entity fp_log_log_24_t1_clk is
  port ( a   : in  std_logic_vector(7 downto 0);
         b   : in  std_logic_vector(15 downto 0);
         r   : out std_logic_vector(28 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_24_t1_clk is
  signal sign_0 : std_logic;
  signal b0_0   : std_logic_vector(14 downto 0);
  signal s_0    : std_logic_vector(15 downto 0);
  component fp_log_log_24_t1_pow is
    port ( x : in  std_logic_vector(14 downto 0);
           r : out std_logic_vector(15 downto 0) );
  end component;

  signal a_1_0    : std_logic_vector(7 downto 0);
  signal sign_1_0 : std_logic;
  signal sgn_1_0  : std_logic;
  signal sgn_1_1  : std_logic;
  signal sgn_1_2  : std_logic;
  signal sgn_1_3  : std_logic;
  signal s_1_0    : std_logic_vector(15 downto 0);
  signal s_1_1    : std_logic_vector(15 downto 0);
  signal k_1_0    : std_logic_vector(20 downto 0);
  signal k_1_1    : std_logic_vector(20 downto 0);
  signal r0_1_3   : std_logic_vector(36 downto 0);
  signal r1_1_3   : std_logic_vector(37 downto 0);
  signal r_1_3    : std_logic_vector(28 downto 0);
  component fp_log_log_24_t1_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(20 downto 0) );
  end component;
begin
  sign_0 <= not b(15);
  b0_0 <= b(14 downto 0) xor (14 downto 0 => sign_0);

  pow : fp_log_log_24_t1_pow
    port map ( x => b0_0,
               r => s_0 );

  a_1_0 <= a(7 downto 0);
  sign_1_0 <= not s_0(15);
  sgn_1_0 <= sign_0 xor sign_1_0;
  s_1_0 <= (s_0(14 downto 0) xor (14 downto 0 => sign_1_0)) & "1";
  t_1 : fp_log_log_24_t1_t1
    port map ( a => a_1_0,
               r => k_1_0 );

  mult_r0_1 : mult_clk
    generic map ( wX    => 21,
                  wY    => 16,
                  first => 0,
                  steps => 2 )
    port map ( nX  => k_1_1,
               nY  => s_1_1,
               nR  => r0_1_3,
               clk => clk );
  
  r1_1_3 <= "0" & r0_1_3;

  r_1_3(20 downto 0) <=
    r1_1_3(37 downto 17) xor (37 downto 17 => (not (sgn_1_3)));
  r_1_3(28 downto 21) <= (28 downto 21 => (not (sgn_1_3)));

  process(clk)
  begin
    if clk'event and clk = '1' then
      s_1_1   <= s_1_0;
      k_1_1   <= k_1_0;
      sgn_1_1 <= sgn_1_0;

      sgn_1_2 <= sgn_1_1;

      sgn_1_3 <= sgn_1_2;
    end if;
  end process;

  r <= r_1_3;
end architecture;


--------------------------------------------------------------------------------
-- PowerAdHoc instance for order-2 powering unit.
-- Decomposition:
--   beta_2 = 12; mu_2 = 18; lambda_2 = 9.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t2_pow is
  port ( x : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of fp_log_log_24_t2_pow is
  signal pp0 : std_logic_vector(16 downto 0);
  signal pp1 : std_logic_vector(16 downto 0);
  signal pp2 : std_logic_vector(16 downto 0);
  signal pp3 : std_logic_vector(16 downto 0);
  signal pp4 : std_logic_vector(16 downto 0);
  signal pp5 : std_logic_vector(16 downto 0);
  signal pp6 : std_logic_vector(16 downto 0);
  signal r0 : std_logic_vector(16 downto 0);
begin
  pp0(16) <= '0';
  pp1(16) <= '0';
  pp2(16) <= '0';
  pp3(16) <= '0';
  pp4(16) <= '0';
  pp5(16) <= '0';
  pp6(16) <= '0';

  pp0(15) <= x(9) and x(10);
  pp1(15) <= x(10);
  pp2(15) <= '0';
  pp3(15) <= '0';
  pp4(15) <= '0';
  pp5(15) <= '0';
  pp6(15) <= '0';

  pp0(14) <= x(8) and x(10);
  pp1(14) <= '0';
  pp2(14) <= '0';
  pp3(14) <= '0';
  pp4(14) <= '0';
  pp5(14) <= '0';
  pp6(14) <= '0';

  pp0(13) <= x(7) and x(10);
  pp1(13) <= x(8) and x(9);
  pp2(13) <= x(9);
  pp3(13) <= '0';
  pp4(13) <= '0';
  pp5(13) <= '0';
  pp6(13) <= '0';

  pp0(12) <= x(6) and x(10);
  pp1(12) <= x(7) and x(9);
  pp2(12) <= '0';
  pp3(12) <= '0';
  pp4(12) <= '0';
  pp5(12) <= '0';
  pp6(12) <= '0';

  pp0(11) <= x(5) and x(10);
  pp1(11) <= x(6) and x(9);
  pp2(11) <= x(7) and x(8);
  pp3(11) <= x(8);
  pp4(11) <= '0';
  pp5(11) <= '0';
  pp6(11) <= '0';

  pp0(10) <= x(4) and x(10);
  pp1(10) <= x(5) and x(9);
  pp2(10) <= x(6) and x(8);
  pp3(10) <= '0';
  pp4(10) <= '0';
  pp5(10) <= '0';
  pp6(10) <= '0';

  pp0(9) <= x(3) and x(10);
  pp1(9) <= x(4) and x(9);
  pp2(9) <= x(5) and x(8);
  pp3(9) <= x(6) and x(7);
  pp4(9) <= x(7);
  pp5(9) <= '0';
  pp6(9) <= '0';

  pp0(8) <= x(2) and x(10);
  pp1(8) <= x(3) and x(9);
  pp2(8) <= x(4) and x(8);
  pp3(8) <= x(5) and x(7);
  pp4(8) <= '0';
  pp5(8) <= '0';
  pp6(8) <= '0';

  pp0(7) <= x(1) and x(10);
  pp1(7) <= x(2) and x(9);
  pp2(7) <= x(3) and x(8);
  pp3(7) <= x(4) and x(7);
  pp4(7) <= x(5) and x(6);
  pp5(7) <= x(6);
  pp6(7) <= '0';

  pp0(6) <= x(0) and x(10);
  pp1(6) <= x(1) and x(9);
  pp2(6) <= x(2) and x(8);
  pp3(6) <= x(3) and x(7);
  pp4(6) <= x(4) and x(6);
  pp5(6) <= '0';
  pp6(6) <= '0';

  pp0(5) <= x(0) and x(9);
  pp1(5) <= x(1) and x(8);
  pp2(5) <= x(2) and x(7);
  pp3(5) <= x(3) and x(6);
  pp4(5) <= x(4) and x(5);
  pp5(5) <= x(5);
  pp6(5) <= x(10);

  pp0(4) <= x(0) and x(8);
  pp1(4) <= x(1) and x(7);
  pp2(4) <= x(2) and x(6);
  pp3(4) <= x(3) and x(5);
  pp4(4) <= x(9);
  pp5(4) <= '0';
  pp6(4) <= '0';

  pp0(3) <= x(0) and x(7);
  pp1(3) <= x(1) and x(6);
  pp2(3) <= x(2) and x(5);
  pp3(3) <= x(3) and x(4);
  pp4(3) <= x(4);
  pp5(3) <= x(8);
  pp6(3) <= '0';

  pp0(2) <= x(0) and x(6);
  pp1(2) <= x(1) and x(5);
  pp2(2) <= x(2) and x(4);
  pp3(2) <= x(7);
  pp4(2) <= '0';
  pp5(2) <= '0';
  pp6(2) <= '0';

  pp0(1) <= x(0) and x(5);
  pp1(1) <= x(1) and x(4);
  pp2(1) <= x(2) and x(3);
  pp3(1) <= x(3);
  pp4(1) <= x(6);
  pp5(1) <= '0';
  pp6(1) <= '0';

  pp0(0) <= x(0) and x(4);
  pp1(0) <= x(1) and x(3);
  pp2(0) <= x(5);
  pp3(0) <= '0';
  pp4(0) <= '0';
  pp5(0) <= '0';
  pp6(0) <= '0';

  r0 <= pp0 + pp1 + pp2 + pp3 + pp4 + pp5 + pp6;
  r <= "1" & r0(16 downto 9);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t2_pow_clk is
  port ( x   : in  std_logic_vector(10 downto 0);
         r   : out std_logic_vector(8 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_24_t2_pow_clk is
  signal pp0 : std_logic_vector(16 downto 0);
  signal pp1 : std_logic_vector(16 downto 0);
  signal pp2 : std_logic_vector(16 downto 0);
  signal pp3 : std_logic_vector(16 downto 0);
  signal pp4 : std_logic_vector(16 downto 0);
  signal pp5 : std_logic_vector(16 downto 0);
  signal pp6 : std_logic_vector(16 downto 0);
  
  signal pp0_0 : std_logic_vector(16 downto 0);
  signal pp0_1 : std_logic_vector(16 downto 0);
  signal pp2_0 : std_logic_vector(16 downto 0);
  signal pp2_1 : std_logic_vector(16 downto 0);
  signal pp4_0 : std_logic_vector(16 downto 0);
  signal pp4_1 : std_logic_vector(16 downto 0);
  signal pp6_0 : std_logic_vector(16 downto 0);
  signal pp6_1 : std_logic_vector(16 downto 0);
  
  signal r0_1 : std_logic_vector(16 downto 0);
begin
  pp0(16) <= '0';
  pp1(16) <= '0';
  pp2(16) <= '0';
  pp3(16) <= '0';
  pp4(16) <= '0';
  pp5(16) <= '0';
  pp6(16) <= '0';

  pp0(15) <= x(9) and x(10);
  pp1(15) <= x(10);
  pp2(15) <= '0';
  pp3(15) <= '0';
  pp4(15) <= '0';
  pp5(15) <= '0';
  pp6(15) <= '0';

  pp0(14) <= x(8) and x(10);
  pp1(14) <= '0';
  pp2(14) <= '0';
  pp3(14) <= '0';
  pp4(14) <= '0';
  pp5(14) <= '0';
  pp6(14) <= '0';

  pp0(13) <= x(7) and x(10);
  pp1(13) <= x(8) and x(9);
  pp2(13) <= x(9);
  pp3(13) <= '0';
  pp4(13) <= '0';
  pp5(13) <= '0';
  pp6(13) <= '0';

  pp0(12) <= x(6) and x(10);
  pp1(12) <= x(7) and x(9);
  pp2(12) <= '0';
  pp3(12) <= '0';
  pp4(12) <= '0';
  pp5(12) <= '0';
  pp6(12) <= '0';

  pp0(11) <= x(5) and x(10);
  pp1(11) <= x(6) and x(9);
  pp2(11) <= x(7) and x(8);
  pp3(11) <= x(8);
  pp4(11) <= '0';
  pp5(11) <= '0';
  pp6(11) <= '0';

  pp0(10) <= x(4) and x(10);
  pp1(10) <= x(5) and x(9);
  pp2(10) <= x(6) and x(8);
  pp3(10) <= '0';
  pp4(10) <= '0';
  pp5(10) <= '0';
  pp6(10) <= '0';

  pp0(9) <= x(3) and x(10);
  pp1(9) <= x(4) and x(9);
  pp2(9) <= x(5) and x(8);
  pp3(9) <= x(6) and x(7);
  pp4(9) <= x(7);
  pp5(9) <= '0';
  pp6(9) <= '0';

  pp0(8) <= x(2) and x(10);
  pp1(8) <= x(3) and x(9);
  pp2(8) <= x(4) and x(8);
  pp3(8) <= x(5) and x(7);
  pp4(8) <= '0';
  pp5(8) <= '0';
  pp6(8) <= '0';

  pp0(7) <= x(1) and x(10);
  pp1(7) <= x(2) and x(9);
  pp2(7) <= x(3) and x(8);
  pp3(7) <= x(4) and x(7);
  pp4(7) <= x(5) and x(6);
  pp5(7) <= x(6);
  pp6(7) <= '0';

  pp0(6) <= x(0) and x(10);
  pp1(6) <= x(1) and x(9);
  pp2(6) <= x(2) and x(8);
  pp3(6) <= x(3) and x(7);
  pp4(6) <= x(4) and x(6);
  pp5(6) <= '0';
  pp6(6) <= '0';

  pp0(5) <= x(0) and x(9);
  pp1(5) <= x(1) and x(8);
  pp2(5) <= x(2) and x(7);
  pp3(5) <= x(3) and x(6);
  pp4(5) <= x(4) and x(5);
  pp5(5) <= x(5);
  pp6(5) <= x(10);

  pp0(4) <= x(0) and x(8);
  pp1(4) <= x(1) and x(7);
  pp2(4) <= x(2) and x(6);
  pp3(4) <= x(3) and x(5);
  pp4(4) <= x(9);
  pp5(4) <= '0';
  pp6(4) <= '0';

  pp0(3) <= x(0) and x(7);
  pp1(3) <= x(1) and x(6);
  pp2(3) <= x(2) and x(5);
  pp3(3) <= x(3) and x(4);
  pp4(3) <= x(4);
  pp5(3) <= x(8);
  pp6(3) <= '0';

  pp0(2) <= x(0) and x(6);
  pp1(2) <= x(1) and x(5);
  pp2(2) <= x(2) and x(4);
  pp3(2) <= x(7);
  pp4(2) <= '0';
  pp5(2) <= '0';
  pp6(2) <= '0';

  pp0(1) <= x(0) and x(5);
  pp1(1) <= x(1) and x(4);
  pp2(1) <= x(2) and x(3);
  pp3(1) <= x(3);
  pp4(1) <= x(6);
  pp5(1) <= '0';
  pp6(1) <= '0';

  pp0(0) <= x(0) and x(4);
  pp1(0) <= x(1) and x(3);
  pp2(0) <= x(5);
  pp3(0) <= '0';
  pp4(0) <= '0';
  pp5(0) <= '0';
  pp6(0) <= '0';

  pp0_0 <= pp0 + pp1;
  pp2_0 <= pp2 + pp3;
  pp4_0 <= pp4 + pp5;
  pp6_0 <= pp6;

  process(clk)
  begin
    if clk'event and clk = '1' then
      pp0_1 <= pp0_0;
      pp2_1 <= pp2_0;
      pp4_1 <= pp4_0;
      pp6_1 <= pp6_0;
    end if;
  end process;
  
  r0_1 <= pp0_1 + pp2_1 + pp4_1 + pp6_1;
  r <= "1" & r0_1(16 downto 9);
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult::Table instance for order-2 term Q_1.
-- Decomposition:
--   alpha_2,1 = 8; wO_2,1 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t2_t1 is
  port ( a : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of fp_log_log_24_t2_t1 is
  signal x : std_logic_vector(7 downto 0);
begin
  x <= a;

  with x select
    r <= "110001000010" when "00000000", -- t[0] = 3138
         "110000001101" when "00000001", -- t[1] = 3085
         "101111011010" when "00000010", -- t[2] = 3034
         "101110101000" when "00000011", -- t[3] = 2984
         "101101110111" when "00000100", -- t[4] = 2935
         "101101000111" when "00000101", -- t[5] = 2887
         "101100011001" when "00000110", -- t[6] = 2841
         "101011101011" when "00000111", -- t[7] = 2795
         "101010111111" when "00001000", -- t[8] = 2751
         "101010010011" when "00001001", -- t[9] = 2707
         "101001101001" when "00001010", -- t[10] = 2665
         "101000111111" when "00001011", -- t[11] = 2623
         "101000010110" when "00001100", -- t[12] = 2582
         "100111101111" when "00001101", -- t[13] = 2543
         "100111001000" when "00001110", -- t[14] = 2504
         "100110100010" when "00001111", -- t[15] = 2466
         "100101111101" when "00010000", -- t[16] = 2429
         "100101011000" when "00010001", -- t[17] = 2392
         "100100110101" when "00010010", -- t[18] = 2357
         "100100010010" when "00010011", -- t[19] = 2322
         "100011110000" when "00010100", -- t[20] = 2288
         "100011001110" when "00010101", -- t[21] = 2254
         "100010101101" when "00010110", -- t[22] = 2221
         "100010001101" when "00010111", -- t[23] = 2189
         "100001101110" when "00011000", -- t[24] = 2158
         "100001001111" when "00011001", -- t[25] = 2127
         "100000110001" when "00011010", -- t[26] = 2097
         "100000010100" when "00011011", -- t[27] = 2068
         "011111110111" when "00011100", -- t[28] = 2039
         "011111011010" when "00011101", -- t[29] = 2010
         "011110111111" when "00011110", -- t[30] = 1983
         "011110100011" when "00011111", -- t[31] = 1955
         "011110001001" when "00100000", -- t[32] = 1929
         "011101101111" when "00100001", -- t[33] = 1903
         "011101010101" when "00100010", -- t[34] = 1877
         "011100111100" when "00100011", -- t[35] = 1852
         "011100100011" when "00100100", -- t[36] = 1827
         "011100001011" when "00100101", -- t[37] = 1803
         "011011110011" when "00100110", -- t[38] = 1779
         "011011011100" when "00100111", -- t[39] = 1756
         "011011000101" when "00101000", -- t[40] = 1733
         "011010101110" when "00101001", -- t[41] = 1710
         "011010011000" when "00101010", -- t[42] = 1688
         "011010000011" when "00101011", -- t[43] = 1667
         "011001101101" when "00101100", -- t[44] = 1645
         "011001011000" when "00101101", -- t[45] = 1624
         "011001000100" when "00101110", -- t[46] = 1604
         "011000110000" when "00101111", -- t[47] = 1584
         "011000011100" when "00110000", -- t[48] = 1564
         "011000001001" when "00110001", -- t[49] = 1545
         "010111110110" when "00110010", -- t[50] = 1526
         "010111100011" when "00110011", -- t[51] = 1507
         "010111010001" when "00110100", -- t[52] = 1489
         "010110111110" when "00110101", -- t[53] = 1470
         "010110101101" when "00110110", -- t[54] = 1453
         "010110011011" when "00110111", -- t[55] = 1435
         "010110001010" when "00111000", -- t[56] = 1418
         "010101111001" when "00111001", -- t[57] = 1401
         "010101101001" when "00111010", -- t[58] = 1385
         "010101011000" when "00111011", -- t[59] = 1368
         "010101001000" when "00111100", -- t[60] = 1352
         "010100111000" when "00111101", -- t[61] = 1336
         "010100101001" when "00111110", -- t[62] = 1321
         "010100011010" when "00111111", -- t[63] = 1306
         "010100001011" when "01000000", -- t[64] = 1291
         "010011111100" when "01000001", -- t[65] = 1276
         "010011101101" when "01000010", -- t[66] = 1261
         "010011011111" when "01000011", -- t[67] = 1247
         "010011010001" when "01000100", -- t[68] = 1233
         "010011000011" when "01000101", -- t[69] = 1219
         "010010110110" when "01000110", -- t[70] = 1206
         "010010101000" when "01000111", -- t[71] = 1192
         "010010011011" when "01001000", -- t[72] = 1179
         "010010001110" when "01001001", -- t[73] = 1166
         "010010000001" when "01001010", -- t[74] = 1153
         "010001110101" when "01001011", -- t[75] = 1141
         "010001101000" when "01001100", -- t[76] = 1128
         "010001011100" when "01001101", -- t[77] = 1116
         "010001010000" when "01001110", -- t[78] = 1104
         "010001000100" when "01001111", -- t[79] = 1092
         "010000111001" when "01010000", -- t[80] = 1081
         "010000101101" when "01010001", -- t[81] = 1069
         "010000100010" when "01010010", -- t[82] = 1058
         "010000010111" when "01010011", -- t[83] = 1047
         "010000001100" when "01010100", -- t[84] = 1036
         "010000000001" when "01010101", -- t[85] = 1025
         "001111110111" when "01010110", -- t[86] = 1015
         "001111101100" when "01010111", -- t[87] = 1004
         "001111100010" when "01011000", -- t[88] = 994
         "001111011000" when "01011001", -- t[89] = 984
         "001111001110" when "01011010", -- t[90] = 974
         "001111000100" when "01011011", -- t[91] = 964
         "001110111010" when "01011100", -- t[92] = 954
         "001110110000" when "01011101", -- t[93] = 944
         "001110100111" when "01011110", -- t[94] = 935
         "001110011110" when "01011111", -- t[95] = 926
         "001110010100" when "01100000", -- t[96] = 916
         "001110001011" when "01100001", -- t[97] = 907
         "001110000010" when "01100010", -- t[98] = 898
         "001101111010" when "01100011", -- t[99] = 890
         "001101110001" when "01100100", -- t[100] = 881
         "001101101000" when "01100101", -- t[101] = 872
         "001101100000" when "01100110", -- t[102] = 864
         "001101011000" when "01100111", -- t[103] = 856
         "001101001111" when "01101000", -- t[104] = 847
         "001101000111" when "01101001", -- t[105] = 839
         "001100111111" when "01101010", -- t[106] = 831
         "001100110111" when "01101011", -- t[107] = 823
         "001100110000" when "01101100", -- t[108] = 816
         "001100101000" when "01101101", -- t[109] = 808
         "001100100000" when "01101110", -- t[110] = 800
         "001100011001" when "01101111", -- t[111] = 793
         "001100010001" when "01110000", -- t[112] = 785
         "001100001010" when "01110001", -- t[113] = 778
         "001100000011" when "01110010", -- t[114] = 771
         "001011111100" when "01110011", -- t[115] = 764
         "001011110101" when "01110100", -- t[116] = 757
         "001011101110" when "01110101", -- t[117] = 750
         "001011100111" when "01110110", -- t[118] = 743
         "001011100001" when "01110111", -- t[119] = 737
         "001011011010" when "01111000", -- t[120] = 730
         "001011010011" when "01111001", -- t[121] = 723
         "001011001101" when "01111010", -- t[122] = 717
         "001011000110" when "01111011", -- t[123] = 710
         "001011000000" when "01111100", -- t[124] = 704
         "001010111010" when "01111101", -- t[125] = 698
         "001010110100" when "01111110", -- t[126] = 692
         "001010101110" when "01111111", -- t[127] = 686
         "001010101000" when "10000000", -- t[128] = 680
         "001010100010" when "10000001", -- t[129] = 674
         "001010011100" when "10000010", -- t[130] = 668
         "001010010110" when "10000011", -- t[131] = 662
         "001010010000" when "10000100", -- t[132] = 656
         "001010001011" when "10000101", -- t[133] = 651
         "001010000101" when "10000110", -- t[134] = 645
         "001010000000" when "10000111", -- t[135] = 640
         "001001111010" when "10001000", -- t[136] = 634
         "001001110101" when "10001001", -- t[137] = 629
         "001001110000" when "10001010", -- t[138] = 624
         "001001101010" when "10001011", -- t[139] = 618
         "001001100101" when "10001100", -- t[140] = 613
         "001001100000" when "10001101", -- t[141] = 608
         "001001011011" when "10001110", -- t[142] = 603
         "001001010110" when "10001111", -- t[143] = 598
         "001001010001" when "10010000", -- t[144] = 593
         "001001001100" when "10010001", -- t[145] = 588
         "001001000111" when "10010010", -- t[146] = 583
         "001001000011" when "10010011", -- t[147] = 579
         "001000111110" when "10010100", -- t[148] = 574
         "001000111001" when "10010101", -- t[149] = 569
         "001000110101" when "10010110", -- t[150] = 565
         "001000110000" when "10010111", -- t[151] = 560
         "001000101100" when "10011000", -- t[152] = 556
         "001000100111" when "10011001", -- t[153] = 551
         "001000100011" when "10011010", -- t[154] = 547
         "001000011110" when "10011011", -- t[155] = 542
         "001000011010" when "10011100", -- t[156] = 538
         "001000010110" when "10011101", -- t[157] = 534
         "001000010010" when "10011110", -- t[158] = 530
         "001000001101" when "10011111", -- t[159] = 525
         "001000001001" when "10100000", -- t[160] = 521
         "001000000101" when "10100001", -- t[161] = 517
         "001000000001" when "10100010", -- t[162] = 513
         "000111111101" when "10100011", -- t[163] = 509
         "000111111001" when "10100100", -- t[164] = 505
         "000111110101" when "10100101", -- t[165] = 501
         "000111110010" when "10100110", -- t[166] = 498
         "000111101110" when "10100111", -- t[167] = 494
         "000111101010" when "10101000", -- t[168] = 490
         "000111100110" when "10101001", -- t[169] = 486
         "000111100011" when "10101010", -- t[170] = 483
         "000111011111" when "10101011", -- t[171] = 479
         "000111011011" when "10101100", -- t[172] = 475
         "000111011000" when "10101101", -- t[173] = 472
         "000111010100" when "10101110", -- t[174] = 468
         "000111010001" when "10101111", -- t[175] = 465
         "000111001101" when "10110000", -- t[176] = 461
         "000111001010" when "10110001", -- t[177] = 458
         "000111000110" when "10110010", -- t[178] = 454
         "000111000011" when "10110011", -- t[179] = 451
         "000111000000" when "10110100", -- t[180] = 448
         "000110111101" when "10110101", -- t[181] = 445
         "000110111001" when "10110110", -- t[182] = 441
         "000110110110" when "10110111", -- t[183] = 438
         "000110110011" when "10111000", -- t[184] = 435
         "000110110000" when "10111001", -- t[185] = 432
         "000110101101" when "10111010", -- t[186] = 429
         "000110101010" when "10111011", -- t[187] = 426
         "000110100110" when "10111100", -- t[188] = 422
         "000110100011" when "10111101", -- t[189] = 419
         "000110100000" when "10111110", -- t[190] = 416
         "000110011110" when "10111111", -- t[191] = 414
         "000110011011" when "11000000", -- t[192] = 411
         "000110011000" when "11000001", -- t[193] = 408
         "000110010101" when "11000010", -- t[194] = 405
         "000110010010" when "11000011", -- t[195] = 402
         "000110001111" when "11000100", -- t[196] = 399
         "000110001100" when "11000101", -- t[197] = 396
         "000110001010" when "11000110", -- t[198] = 394
         "000110000111" when "11000111", -- t[199] = 391
         "000110000100" when "11001000", -- t[200] = 388
         "000110000001" when "11001001", -- t[201] = 385
         "000101111111" when "11001010", -- t[202] = 383
         "000101111100" when "11001011", -- t[203] = 380
         "000101111010" when "11001100", -- t[204] = 378
         "000101110111" when "11001101", -- t[205] = 375
         "000101110100" when "11001110", -- t[206] = 372
         "000101110010" when "11001111", -- t[207] = 370
         "000101101111" when "11010000", -- t[208] = 367
         "000101101101" when "11010001", -- t[209] = 365
         "000101101011" when "11010010", -- t[210] = 363
         "000101101000" when "11010011", -- t[211] = 360
         "000101100110" when "11010100", -- t[212] = 358
         "000101100011" when "11010101", -- t[213] = 355
         "000101100001" when "11010110", -- t[214] = 353
         "000101011111" when "11010111", -- t[215] = 351
         "000101011100" when "11011000", -- t[216] = 348
         "000101011010" when "11011001", -- t[217] = 346
         "000101011000" when "11011010", -- t[218] = 344
         "000101010101" when "11011011", -- t[219] = 341
         "000101010011" when "11011100", -- t[220] = 339
         "000101010001" when "11011101", -- t[221] = 337
         "000101001111" when "11011110", -- t[222] = 335
         "000101001101" when "11011111", -- t[223] = 333
         "000101001010" when "11100000", -- t[224] = 330
         "000101001000" when "11100001", -- t[225] = 328
         "000101000110" when "11100010", -- t[226] = 326
         "000101000100" when "11100011", -- t[227] = 324
         "000101000010" when "11100100", -- t[228] = 322
         "000101000000" when "11100101", -- t[229] = 320
         "000100111110" when "11100110", -- t[230] = 318
         "000100111100" when "11100111", -- t[231] = 316
         "000100111010" when "11101000", -- t[232] = 314
         "000100111000" when "11101001", -- t[233] = 312
         "000100110110" when "11101010", -- t[234] = 310
         "000100110100" when "11101011", -- t[235] = 308
         "000100110010" when "11101100", -- t[236] = 306
         "000100110000" when "11101101", -- t[237] = 304
         "000100101110" when "11101110", -- t[238] = 302
         "000100101100" when "11101111", -- t[239] = 300
         "000100101011" when "11110000", -- t[240] = 299
         "000100101001" when "11110001", -- t[241] = 297
         "000100100111" when "11110010", -- t[242] = 295
         "000100100101" when "11110011", -- t[243] = 293
         "000100100011" when "11110100", -- t[244] = 291
         "000100100001" when "11110101", -- t[245] = 289
         "000100100000" when "11110110", -- t[246] = 288
         "000100011110" when "11110111", -- t[247] = 286
         "000100011100" when "11111000", -- t[248] = 284
         "000100011010" when "11111001", -- t[249] = 282
         "000100011001" when "11111010", -- t[250] = 281
         "000100010111" when "11111011", -- t[251] = 279
         "000100010101" when "11111100", -- t[252] = 277
         "000100010100" when "11111101", -- t[253] = 276
         "000100010010" when "11111110", -- t[254] = 274
         "000100010000" when "11111111", -- t[255] = 272
         "------------" when others;
end architecture;


--------------------------------------------------------------------------------
-- TermPowMult instance for order-2 term.
-- Decomposition:
--   alpha_2 = 8; beta_2 = 12; lambda_2 = 9;  m_2 = 1;
--   Pow   (AdHoc);
--   Q_2,1 (Mult): alpha_2,1 = 8; rho_2,1 = 0; sigma_2,1 = 9; wO_2,1 = 12.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t2 is
  port ( a : in  std_logic_vector(7 downto 0);
         b : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(28 downto 0) );
end entity;

architecture arch of fp_log_log_24_t2 is
  signal sign   : std_logic;
  signal b0     : std_logic_vector(10 downto 0);
  signal s      : std_logic_vector(8 downto 0);
  component fp_log_log_24_t2_pow is
    port ( x : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  signal a_1    : std_logic_vector(7 downto 0);
  signal sign_1 : std_logic;
  signal s_1    : std_logic_vector(7 downto 0);
  signal k_1    : std_logic_vector(11 downto 0);
  signal r0_1   : std_logic_vector(21 downto 0);
  signal r_1    : std_logic_vector(28 downto 0);
  component fp_log_log_24_t2_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;
begin
  sign <= not b(11);
  b0 <= b(10 downto 0) xor (10 downto 0 => sign);

  pow : fp_log_log_24_t2_pow
    port map ( x => b0,
               r => s );

  a_1 <= a(7 downto 0);
  sign_1 <= not s(8);
  s_1 <= s(7 downto 0) xor (7 downto 0 => sign_1);
  t_1 : fp_log_log_24_t2_t1
    port map ( a => a_1,
               r => k_1 );
  r0_1 <= "0" & (k_1 * (s_1 & "1"));
  r_1(11 downto 0) <=
    r0_1(21 downto 10) xor (21 downto 10 => ((sign_1)));
  r_1(28 downto 12) <= (28 downto 12 => ((sign_1)));

  r <= r_1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_fp_log.all;

entity fp_log_log_24_t2_clk is
  port ( a   : in  std_logic_vector(7 downto 0);
         b   : in  std_logic_vector(11 downto 0);
         r   : out std_logic_vector(28 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_24_t2_clk is
  signal sign_0 : std_logic;
  signal b0_0   : std_logic_vector(10 downto 0);
  signal s_1    : std_logic_vector(8 downto 0);
  component fp_log_log_24_t2_pow_clk is
    port ( x   : in  std_logic_vector(10 downto 0);
           r   : out std_logic_vector(8 downto 0);
           clk : in  std_logic );
  end component;

  signal a_1_0    : std_logic_vector(7 downto 0);
  signal a_1_1    : std_logic_vector(7 downto 0);
  signal sign_1_1 : std_logic;
  signal sign_1_2 : std_logic;
  signal sign_1_3 : std_logic;
  signal sign_1_4 : std_logic;
  signal s_1_1    : std_logic_vector(8 downto 0);
  signal s_1_2    : std_logic_vector(8 downto 0);
  signal k_1_1    : std_logic_vector(11 downto 0);
  signal k_1_2    : std_logic_vector(11 downto 0);
  signal r0_1_4   : std_logic_vector(20 downto 0);
  signal r1_1_4   : std_logic_vector(21 downto 0);
  signal r_1_4    : std_logic_vector(28 downto 0);
  component fp_log_log_24_t2_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;
begin
  sign_0 <= not b(11);
  b0_0 <= b(10 downto 0) xor (10 downto 0 => sign_0);

  pow : fp_log_log_24_t2_pow_clk
    port map ( x   => b0_0,
               r   => s_1,
               clk => clk );

  a_1_0 <= a(7 downto 0);
  sign_1_1 <= not s_1(8);
  s_1_1 <= (s_1(7 downto 0) xor (7 downto 0 => sign_1_1)) & "1";
  t_1 : fp_log_log_24_t2_t1
    port map ( a => a_1_1,
               r => k_1_1 );

  mult_r0_1 : mult_clk
    generic map ( wX    => 12,
                  wY    => 9,
                  first => 0,
                  steps => 2 )
    port map ( nX  => k_1_2,
               nY  => s_1_2,
               nR  => r0_1_4,
               clk => clk );
  
  r1_1_4 <= "0" & r0_1_4;

  r_1_4(11 downto 0) <=
    r1_1_4(21 downto 10) xor (21 downto 10 => ((sign_1_4)));
  r_1_4(28 downto 12) <= (28 downto 12 => ((sign_1_4)));

  process(clk)
  begin
    if clk'event and clk = '1' then
      a_1_1    <= a_1_0;
      
      sign_1_2 <= sign_1_1;
      s_1_2    <= s_1_1;
      k_1_2    <= k_1_1;

      sign_1_3 <= sign_1_2;

      sign_1_4 <= sign_1_3;
    end if;
  end process;

  r <= r_1_4;
end architecture;


--------------------------------------------------------------------------------
-- TermROM instance for order-3 term.
-- Decomposition:
--   alpha_3 = 2; beta_3 = 3 (1+2); wO_3 = 2.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_t3 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(28 downto 0) );
end entity;

architecture arch of fp_log_log_24_t3 is
  signal sign : std_logic;
  signal b0   : std_logic_vector(1 downto 0);
  signal x0   : std_logic_vector(3 downto 0);
  signal r0   : std_logic_vector(1 downto 0);
begin
  sign <= not b(2);
  b0 <= b(1 downto 0) xor (1 downto 0 => sign);
  x0 <= a & b0;

  with x0 select
    r0 <= "11" when "0000", -- t[0] = -1
          "11" when "0001", -- t[1] = -1
          "11" when "0010", -- t[2] = -1
          "01" when "0011", -- t[3] = -3
          "11" when "0100", -- t[4] = -1
          "11" when "0101", -- t[5] = -1
          "11" when "0110", -- t[6] = -1
          "11" when "0111", -- t[7] = -1
          "11" when "1000", -- t[8] = -1
          "11" when "1001", -- t[9] = -1
          "11" when "1010", -- t[10] = -1
          "11" when "1011", -- t[11] = -1
          "11" when "1100", -- t[12] = -1
          "11" when "1101", -- t[13] = -1
          "11" when "1110", -- t[14] = -1
          "11" when "1111", -- t[15] = -1
          "--" when others;

  r(1 downto 0) <= r0 xor (1 downto 0 => (not sign));
  r(28 downto 2) <= (28 downto 2 => (not sign));
end architecture;


--------------------------------------------------------------------------------
-- HOTBM main component.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24 is
  port ( x : in  std_logic_vector(23 downto 0);
         r : out std_logic_vector(28 downto 0) );
end entity;

architecture arch of fp_log_log_24 is
  signal a_0 : std_logic_vector(7 downto 0);
  signal r_0 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t0 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(28 downto 0) );
  end component;

  signal a_1 : std_logic_vector(7 downto 0);
  signal b_1 : std_logic_vector(15 downto 0);
  signal r_1 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t1 is
    port ( a : in  std_logic_vector(7 downto 0);
           b : in  std_logic_vector(15 downto 0);
           r : out std_logic_vector(28 downto 0) );
  end component;

  signal a_2 : std_logic_vector(7 downto 0);
  signal b_2 : std_logic_vector(11 downto 0);
  signal r_2 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t2 is
    port ( a : in  std_logic_vector(7 downto 0);
           b : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(28 downto 0) );
  end component;

  signal a_3 : std_logic_vector(1 downto 0);
  signal b_3 : std_logic_vector(2 downto 0);
  signal r_3 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(28 downto 0) );
  end component;

begin
  a_0 <= x(23 downto 16);
  t_0 : fp_log_log_24_t0
    port map ( a => a_0,
               r => r_0 );

  a_1 <= x(23 downto 16);
  b_1 <= x(15 downto 0);
  t_1 : fp_log_log_24_t1
    port map ( a => a_1,
               b => b_1,
               r => r_1 );

  a_2 <= x(23 downto 16);
  b_2 <= x(15 downto 4);
  t_2 : fp_log_log_24_t2
    port map ( a => a_2,
               b => b_2,
               r => r_2 );

  a_3 <= x(23 downto 22);
  b_3 <= x(15 downto 13);
  t_3 : fp_log_log_24_t3
    port map ( a => a_3,
               b => b_3,
               r => r_3 );

  r <= r_0 + r_1 + r_2 + r_3;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fp_log_log_24_clk is
  port ( x   : in  std_logic_vector(23 downto 0);
         r   : out std_logic_vector(28 downto 0);
         clk : in  std_logic );
end entity;

architecture arch of fp_log_log_24_clk is
  signal x_0 : std_logic_vector(23 downto 0);
  signal x_1 : std_logic_vector(23 downto 0);
  signal x_2 : std_logic_vector(23 downto 0);
  signal x_3 : std_logic_vector(23 downto 0);
  signal x_4 : std_logic_vector(23 downto 0);
  
  signal a_0_4 : std_logic_vector(7 downto 0);
  signal r_0_4 : std_logic_vector(28 downto 0);
  signal r_0_5 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t0 is
    port ( a : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(28 downto 0) );
  end component;

  signal a_1_1 : std_logic_vector(7 downto 0);
  signal b_1_1 : std_logic_vector(15 downto 0);
  signal r_1_4 : std_logic_vector(28 downto 0);
  signal r_1_5 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t1_clk is
    port ( a   : in  std_logic_vector(7 downto 0);
           b   : in  std_logic_vector(15 downto 0);
           r   : out std_logic_vector(28 downto 0);
           clk : in  std_logic );
  end component;

  signal a_2_0 : std_logic_vector(7 downto 0);
  signal b_2_0 : std_logic_vector(11 downto 0);
  signal r_2_4 : std_logic_vector(28 downto 0);
  signal r_2_5 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t2_clk is
    port ( a   : in  std_logic_vector(7 downto 0);
           b   : in  std_logic_vector(11 downto 0);
           r   : out std_logic_vector(28 downto 0);
           clk : in  std_logic );
  end component;

  signal a_3_4 : std_logic_vector(1 downto 0);
  signal b_3_4 : std_logic_vector(2 downto 0);
  signal r_3_4 : std_logic_vector(28 downto 0);
  signal r_3_5 : std_logic_vector(28 downto 0);
  component fp_log_log_24_t3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(28 downto 0) );
  end component;

begin
  x_0 <= x;
  
  a_0_4 <= x_4(23 downto 16);
  t_0 : fp_log_log_24_t0
    port map ( a => a_0_4,
               r => r_0_4 );

  a_1_1 <= x_1(23 downto 16);
  b_1_1 <= x_1(15 downto 0);
  t_1 : fp_log_log_24_t1_clk
    port map ( a   => a_1_1,
               b   => b_1_1,
               r   => r_1_4,
               clk => clk );

  a_2_0 <= x_0(23 downto 16);
  b_2_0 <= x_0(15 downto 4);
  t_2 : fp_log_log_24_t2_clk
    port map ( a   => a_2_0,
               b   => b_2_0,
               r   => r_2_4,
               clk => clk );

  a_3_4 <= x_4(23 downto 22);
  b_3_4 <= x_4(15 downto 13);
  t_3 : fp_log_log_24_t3
    port map ( a => a_3_4,
               b => b_3_4,
               r => r_3_4 );

  process(clk)
  begin
    if clk'event and clk = '1' then
      x_1   <= x_0;
      x_2   <= x_1;
      x_3   <= x_2;
      x_4   <= x_3;
      r_0_5 <= r_0_4;
      r_1_5 <= r_1_4;
      r_2_5 <= r_2_4;
      r_3_5 <= r_3_4;
    end if;
  end process;

  r <= r_0_5 + r_1_5 + r_2_5 + r_3_5;
end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_fp_log.all;
use fplib.pkg_fp_log_log.all;

entity fp_log_log is
  generic ( w : positive );
  port ( nX    : in  std_logic_vector(w-1 downto 0);
         nLogX : out std_logic_vector(w+fp_log_log_g(w) downto 0) );
end entity;

architecture arch of fp_log_log is
begin

  log_7 : if w = 7 generate
    log : fp_log_log_7
      port map ( nX    => nX,
                 nLogX => nLogX );
  end generate;

  log_8 : if w = 8 generate
    log : fp_log_log_8
      port map ( nX    => nX,
                 nLogX => nLogX );
  end generate;

  log_9 : if w = 9 generate
    log : fp_log_log_9
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_10 : if w = 10 generate
    log : fp_log_log_10
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_11 : if w = 11 generate
    log : fp_log_log_11
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_12 : if w = 12 generate
    log : fp_log_log_12
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_13 : if w = 13 generate
    log : fp_log_log_13
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_14 : if w = 14 generate
    log : fp_log_log_14
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_15 : if w = 15 generate
    log : fp_log_log_15
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_16 : if w = 16 generate
    log : fp_log_log_16
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_17 : if w = 17 generate
    log : fp_log_log_17
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_18 : if w = 18 generate
    log : fp_log_log_18
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_19 : if w = 19 generate
    log : fp_log_log_19
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_20 : if w = 20 generate
    log : fp_log_log_20
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_21 : if w = 21 generate
    log : fp_log_log_21
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_22 : if w = 22 generate
    log : fp_log_log_22
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_23 : if w = 23 generate
    log : fp_log_log_23
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_24 : if w = 24 generate
    log : fp_log_log_24
      port map ( x => nX,
                 r => nLogX );
  end generate;

end architecture;

-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_fp_log.all;
use fplib.pkg_fp_log_log.all;

entity fp_log_log_clk is
  generic ( w : positive );
  port ( nX    : in  std_logic_vector(w-1 downto 0);
         nLogX : out std_logic_vector(w+fp_log_log_g(w) downto 0);
         clk   : in  std_logic );
end entity;

architecture arch of fp_log_log_clk is
begin

  log_7 : if w = 7 generate
    log : fp_log_log_7
      port map ( nX    => nX,
                 nLogX => nLogX );
  end generate;

  log_8 : if w = 8 generate
    log : fp_log_log_8
      port map ( nX    => nX,
                 nLogX => nLogX );
  end generate;

  log_9 : if w = 9 generate
    log : fp_log_log_9
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_10 : if w = 10 generate
    log : fp_log_log_10
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_11 : if w = 11 generate
    log : fp_log_log_11_clk
      port map ( x   => nX,
                 r   => nLogX,
                 clk => clk );
  end generate;

  log_12 : if w = 12 generate
    log : fp_log_log_12
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_13 : if w = 13 generate
    log : fp_log_log_13
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_14 : if w = 14 generate
    log : fp_log_log_14
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_15 : if w = 15 generate
    log : fp_log_log_15
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_16 : if w = 16 generate
    log : fp_log_log_16
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_17 : if w = 17 generate
    log : fp_log_log_17
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_18 : if w = 18 generate
    log : fp_log_log_18_clk
      port map ( x   => nX,
                 r   => nLogX,
                 clk => clk );
  end generate;

  log_19 : if w = 19 generate
    log : fp_log_log_19
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_20 : if w = 20 generate
    log : fp_log_log_20
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_21 : if w = 21 generate
    log : fp_log_log_21
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_22 : if w = 22 generate
    log : fp_log_log_22
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_23 : if w = 23 generate
    log : fp_log_log_23
      port map ( x => nX,
                 r => nLogX );
  end generate;

  log_24 : if w = 24 generate
    log : fp_log_log_24_clk
      port map ( x   => nX,
                 r   => nLogX,
                 clk => clk );
  end generate;

end architecture;
